// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module BlackBoxRom
#(
    parameter  addrWidth = 11,
               instrWidth = 32
)
(
    input wire [addrWidth-1:0] addressEven,
    input wire [addrWidth-1:0] addressOdd,
    output reg [instrWidth-1:0] instructionEven,
    output reg [instrWidth-1:0] instructionOdd
);
        
always @(*) case (addressEven)
	0: instructionEven = 32'h54;
	1: instructionEven = 32'h20700;
	2: instructionEven = 32'h20800;
	3: instructionEven = 32'h2402025;
	4: instructionEven = 32'h87c20000;
	5: instructionEven = 32'h2821085;
	6: instructionEven = 32'h2021062;
	7: instructionEven = 32'hf0010000;
	8: instructionEven = 32'h80000000;
	9: instructionEven = 32'h400000;
	10: instructionEven = 32'h4000017;
	11: instructionEven = 32'h4ac;
	12: instructionEven = 32'h2520038;
	13: instructionEven = 32'h2c5fd08;
	14: instructionEven = 32'h2c5f481;
	15: instructionEven = 32'h2c5f480;
	16: instructionEven = 32'h2c5fb04;
	17: instructionEven = 32'h2c5fc06;
	18: instructionEven = 32'h87c20000;
	19: instructionEven = 32'h2821083;
	20: instructionEven = 32'h2022081;
	21: instructionEven = 32'hf0020000;
	22: instructionEven = 32'h400000;
	23: instructionEven = 32'h2022062;
	24: instructionEven = 32'h2c60005;
	25: instructionEven = 32'h87c20000;
	26: instructionEven = 32'h2821080;
	27: instructionEven = 32'h2021031;
	28: instructionEven = 32'h87c20000;
	29: instructionEven = 32'h2841080;
	30: instructionEven = 32'hc42004;
	31: instructionEven = 32'h2841080;
	32: instructionEven = 32'hc42004;
	33: instructionEven = 32'h2841080;
	34: instructionEven = 32'hc42004;
	35: instructionEven = 32'h2821080;
	36: instructionEven = 32'hc21004;
	37: instructionEven = 32'h40001;
	38: instructionEven = 32'hf0000000;
	39: instructionEven = 32'h400000;
	40: instructionEven = 32'h2c61109;
	41: instructionEven = 32'h400000;
	42: instructionEven = 32'hcbffff7;
	43: instructionEven = 32'h400000;
	44: instructionEven = 32'hcbffffd;
	45: instructionEven = 32'h87c40000;
	46: instructionEven = 32'h2842082;
	47: instructionEven = 32'h2022060;
	48: instructionEven = 32'h20010;
	49: instructionEven = 32'hc22004;
	50: instructionEven = 32'h460001;
	51: instructionEven = 32'h2c61007;
	52: instructionEven = 32'h20010;
	53: instructionEven = 32'hf0000000;
	54: instructionEven = 32'h42001;
	55: instructionEven = 32'hcbffff4;
	56: instructionEven = 32'h2021031;
	57: instructionEven = 32'h40001;
	58: instructionEven = 32'h4000143;
	59: instructionEven = 32'h87c20000;
	60: instructionEven = 32'h282108c;
	61: instructionEven = 32'h2021264;
	62: instructionEven = 32'hc80000d;
	63: instructionEven = 32'h10000;
	64: instructionEven = 32'h400000;
	65: instructionEven = 32'h87c40000;
	66: instructionEven = 32'h284208c;
	67: instructionEven = 32'h1042002;
	68: instructionEven = 32'hcbffff5;
	69: instructionEven = 32'hf0000000;
	70: instructionEven = 32'h400000;
	71: instructionEven = 32'h4c800008;
	72: instructionEven = 32'hf0000000;
	73: instructionEven = 32'h40002;
	74: instructionEven = 32'hc21004;
	75: instructionEven = 32'h20002;
	76: instructionEven = 32'h87c40000;
	77: instructionEven = 32'h2842082;
	78: instructionEven = 32'h2022164;
	79: instructionEven = 32'hc41004;
	80: instructionEven = 32'h400000;
	81: instructionEven = 32'hcbffffc;
	82: instructionEven = 32'hf0000000;
	83: instructionEven = 32'h21001;
	84: instructionEven = 32'hcbffff6;
	85: instructionEven = 32'h200ff;
	86: instructionEven = 32'hc800023;
	87: instructionEven = 32'hf0010000;
	88: instructionEven = 32'h440001;
	89: instructionEven = 32'hcfc40000;
	90: instructionEven = 32'hcfc20000;
	91: instructionEven = 32'h4ac22085;
	92: instructionEven = 32'h400000;
	93: instructionEven = 32'h400000;
	94: instructionEven = 32'h87c40000;
	95: instructionEven = 32'h2842085;
	96: instructionEven = 32'h2022062;
	97: instructionEven = 32'hf0010000;
	98: instructionEven = 32'h80000000;
	99: instructionEven = 32'h400000;
	100: instructionEven = 32'h87c40000;
	101: instructionEven = 32'h2842080;
	102: instructionEven = 32'hc42004;
	103: instructionEven = 32'h1c210ff;
	104: instructionEven = 32'hf0000000;
	105: instructionEven = 32'h400000;
	106: instructionEven = 32'h4c800012;
	107: instructionEven = 32'h87c20000;
	108: instructionEven = 32'h2821080;
	109: instructionEven = 32'hc21004;
	110: instructionEven = 32'h2820185;
	111: instructionEven = 32'h2021261;
	112: instructionEven = 32'h87c20000;
	113: instructionEven = 32'h2821080;
	114: instructionEven = 32'hc21004;
	115: instructionEven = 32'h87c60000;
	116: instructionEven = 32'h2863082;
	117: instructionEven = 32'h2023164;
	118: instructionEven = 32'hc62004;
	119: instructionEven = 32'h400000;
	120: instructionEven = 32'hc800006;
	121: instructionEven = 32'h2863189;
	122: instructionEven = 32'h2023261;
	123: instructionEven = 32'h87c60000;
	124: instructionEven = 32'h2863082;
	125: instructionEven = 32'h20221b4;
	126: instructionEven = 32'h87c40000;
	127: instructionEven = 32'h2842080;
	128: instructionEven = 32'h2022036;
	129: instructionEven = 32'h87c40000;
	130: instructionEven = 32'h2c22001;
	131: instructionEven = 32'hf0080000;
	132: instructionEven = 32'h400000;
	133: instructionEven = 32'h4cbffffb;
	134: instructionEven = 32'h87c60000;
	135: instructionEven = 32'h2c23101;
	136: instructionEven = 32'hf0080000;
	137: instructionEven = 32'h400000;
	138: instructionEven = 32'h4cbffffb;
	139: instructionEven = 32'hf0080000;
	140: instructionEven = 32'h20004;
	141: instructionEven = 32'h87c40000;
	142: instructionEven = 32'h2842082;
	143: instructionEven = 32'h2022164;
	144: instructionEven = 32'hc41004;
	145: instructionEven = 32'h400000;
	146: instructionEven = 32'hcbffffc;
	147: instructionEven = 32'hf0000000;
	148: instructionEven = 32'h21001;
	149: instructionEven = 32'hcbffff6;
	150: instructionEven = 32'hf0010000;
	151: instructionEven = 32'h4400001;
	152: instructionEven = 32'h20002;
	153: instructionEven = 32'h2adf104;
	154: instructionEven = 32'h2b1f106;
	155: instructionEven = 32'h2b5f108;
	156: instructionEven = 32'h2abf103;
	157: instructionEven = 32'h293f101;
	158: instructionEven = 32'h2409027;
	159: instructionEven = 32'h6400000;
	160: instructionEven = 32'h2409020;
	161: instructionEven = 32'h340;
	162: instructionEven = 32'h2520038;
	163: instructionEven = 32'h87c20000;
	164: instructionEven = 32'h2c41000;
	165: instructionEven = 32'h2520037;
	166: instructionEven = 32'h2520030;
	167: instructionEven = 32'h2c5fa88;
	168: instructionEven = 32'h2c5fb8a;
	169: instructionEven = 32'h2c5fc8c;
	170: instructionEven = 32'h2c5fd8e;
	171: instructionEven = 32'h87c21000;
	172: instructionEven = 32'h40020;
	173: instructionEven = 32'h87c40000;
	174: instructionEven = 32'h2822100;
	175: instructionEven = 32'h21001;
	176: instructionEven = 32'h403be;
	177: instructionEven = 32'hcbffff4;
	178: instructionEven = 32'h20404;
	179: instructionEven = 32'h460001;
	180: instructionEven = 32'h360000;
	181: instructionEven = 32'h2a0000;
	182: instructionEven = 32'h300000;
	183: instructionEven = 32'h2c5f000;
	184: instructionEven = 32'h87c20000;
	185: instructionEven = 32'h2c41000;
	186: instructionEven = 32'h2c5f084;
	187: instructionEven = 32'h20000;
	188: instructionEven = 32'h322000;
	189: instructionEven = 32'h4400214;
	190: instructionEven = 32'hf0090000;
	191: instructionEven = 32'h2c4000;
	192: instructionEven = 32'h203c060;
	193: instructionEven = 32'h80000;
	194: instructionEven = 32'h40003;
	195: instructionEven = 32'hc800005;
	196: instructionEven = 32'h4c0005d;
	197: instructionEven = 32'h59000;
	198: instructionEven = 32'h2022b35;
	199: instructionEven = 32'h2081c82;
	200: instructionEven = 32'h1044001;
	201: instructionEven = 32'h87c42002;
	202: instructionEven = 32'h202104a;
	203: instructionEven = 32'h82000;
	204: instructionEven = 32'h2023031;
	205: instructionEven = 32'hc75003;
	206: instructionEven = 32'h1c63018;
	207: instructionEven = 32'h2021183;
	208: instructionEven = 32'h20004;
	209: instructionEven = 32'hcc00013;
	210: instructionEven = 32'h75001;
	211: instructionEven = 32'hc800013;
	212: instructionEven = 32'h2021db4;
	213: instructionEven = 32'h87c3b00d;
	214: instructionEven = 32'h2861100;
	215: instructionEven = 32'h6003005;
	216: instructionEven = 32'h400000;
	217: instructionEven = 32'h4c00033;
	218: instructionEven = 32'h77000;
	219: instructionEven = 32'h87c21007;
	220: instructionEven = 32'h2c61280;
	221: instructionEven = 32'h283f101;
	222: instructionEven = 32'h85000;
	223: instructionEven = 32'h305000;
	224: instructionEven = 32'h345000;
	225: instructionEven = 32'h400000;
	226: instructionEven = 32'h60000;
	227: instructionEven = 32'h205b2e0;
	228: instructionEven = 32'h4c800015;
	229: instructionEven = 32'h87c63007;
	230: instructionEven = 32'h203a1b5;
	231: instructionEven = 32'h400000;
	232: instructionEven = 32'h2098180;
	233: instructionEven = 32'h2023d34;
	234: instructionEven = 32'h87c84007;
	235: instructionEven = 32'h2c64000;
	236: instructionEven = 32'h2a0000;
	237: instructionEven = 32'h4c00005;
	238: instructionEven = 32'h2c5f180;
	239: instructionEven = 32'h2a3000;
	240: instructionEven = 32'h2023060;
	241: instructionEven = 32'h2c5f283;
	242: instructionEven = 32'h77000;
	243: instructionEven = 32'h20360b1;
	244: instructionEven = 32'h96001;
	245: instructionEven = 32'h87c20000;
	246: instructionEven = 32'h2821080;
	247: instructionEven = 32'h2021036;
	248: instructionEven = 32'h202200b;
	249: instructionEven = 32'h87ca0000;
	250: instructionEven = 32'h20230b1;
	251: instructionEven = 32'h2c25101;
	252: instructionEven = 32'h283f100;
	253: instructionEven = 32'h400000;
	254: instructionEven = 32'hcffff7b;
	255: instructionEven = 32'h43000;
	256: instructionEven = 32'h400000;
	257: instructionEven = 32'h2aff10a;
	258: instructionEven = 32'h2b3f10c;
	259: instructionEven = 32'h2b7f10e;
	260: instructionEven = 32'h293f107;
	261: instructionEven = 32'h2409028;
	262: instructionEven = 32'h400000;
	263: instructionEven = 32'h293f105;
	264: instructionEven = 32'h400000;
	265: instructionEven = 32'h3ff040;
	266: instructionEven = 32'h87c20000;
	267: instructionEven = 32'h87c40000;
	268: instructionEven = 32'h2821100;
	269: instructionEven = 32'h24c0030;
	270: instructionEven = 32'hc800055;
	271: instructionEven = 32'h20408;
	272: instructionEven = 32'h400000;
	273: instructionEven = 32'h2021466;
	274: instructionEven = 32'h400000;
	275: instructionEven = 32'h87c20000;
	276: instructionEven = 32'h2821080;
	277: instructionEven = 32'h1c21002;
	278: instructionEven = 32'hcbffffa;
	279: instructionEven = 32'hf0080000;
	280: instructionEven = 32'h87c40000;
	281: instructionEven = 32'h87c21006;
	282: instructionEven = 32'h2c42080;
	283: instructionEven = 32'h87c20000;
	284: instructionEven = 32'h2821080;
	285: instructionEven = 32'h1c21002;
	286: instructionEven = 32'hcbffffa;
	287: instructionEven = 32'h87c20000;
	288: instructionEven = 32'hcc0000e;
	289: instructionEven = 32'h400000;
	290: instructionEven = 32'h20000;
	291: instructionEven = 32'h400000;
	292: instructionEven = 32'h20004;
	293: instructionEven = 32'h23001;
	294: instructionEven = 32'h1c213ff;
	295: instructionEven = 32'h87c40000;
	296: instructionEven = 32'h2842080;
	297: instructionEven = 32'h1c42002;
	298: instructionEven = 32'hcbffffa;
	299: instructionEven = 32'hf0080000;
	300: instructionEven = 32'h400000;
	301: instructionEven = 32'h1c42300;
	302: instructionEven = 32'h87c40000;
	303: instructionEven = 32'h2842100;
	304: instructionEven = 32'h2063080;
	305: instructionEven = 32'h1c813ff;
	306: instructionEven = 32'h20004;
	307: instructionEven = 32'h87ca2000;
	308: instructionEven = 32'h2d45200;
	309: instructionEven = 32'h21001;
	310: instructionEven = 32'h42001;
	311: instructionEven = 32'h87c20000;
	312: instructionEven = 32'h2c41100;
	313: instructionEven = 32'h20404;
	314: instructionEven = 32'h400000;
	315: instructionEven = 32'h20004;
	316: instructionEven = 32'h1c633ff;
	317: instructionEven = 32'h2821900;
	318: instructionEven = 32'h2406020;
	319: instructionEven = 32'h0;
	320: instructionEven = 32'h0;
	321: instructionEven = 32'h0;
	322: instructionEven = 32'h0;
	323: instructionEven = 32'h0;
	324: instructionEven = 32'h0;
	325: instructionEven = 32'h0;
	326: instructionEven = 32'h0;
	327: instructionEven = 32'h0;
	328: instructionEven = 32'h0;
	329: instructionEven = 32'h0;
	330: instructionEven = 32'h0;
	331: instructionEven = 32'h0;
	332: instructionEven = 32'h0;
	333: instructionEven = 32'h0;
	334: instructionEven = 32'h0;
	335: instructionEven = 32'h0;
	336: instructionEven = 32'h0;
	337: instructionEven = 32'h0;
	338: instructionEven = 32'h0;
	339: instructionEven = 32'h0;
	340: instructionEven = 32'h0;
	341: instructionEven = 32'h0;
	342: instructionEven = 32'h0;
	343: instructionEven = 32'h0;
	344: instructionEven = 32'h0;
	345: instructionEven = 32'h0;
	346: instructionEven = 32'h0;
	347: instructionEven = 32'h0;
	348: instructionEven = 32'h0;
	349: instructionEven = 32'h0;
	350: instructionEven = 32'h0;
	351: instructionEven = 32'h0;
	352: instructionEven = 32'h0;
	353: instructionEven = 32'h0;
	354: instructionEven = 32'h0;
	355: instructionEven = 32'h0;
	356: instructionEven = 32'h0;
	357: instructionEven = 32'h0;
	358: instructionEven = 32'h0;
	359: instructionEven = 32'h0;
	360: instructionEven = 32'h0;
	361: instructionEven = 32'h0;
	362: instructionEven = 32'h0;
	363: instructionEven = 32'h0;
	364: instructionEven = 32'h0;
	365: instructionEven = 32'h0;
	366: instructionEven = 32'h0;
	367: instructionEven = 32'h0;
	368: instructionEven = 32'h0;
	369: instructionEven = 32'h0;
	370: instructionEven = 32'h0;
	371: instructionEven = 32'h0;
	372: instructionEven = 32'h0;
	373: instructionEven = 32'h0;
	374: instructionEven = 32'h0;
	375: instructionEven = 32'h0;
	376: instructionEven = 32'h0;
	377: instructionEven = 32'h0;
	378: instructionEven = 32'h0;
	379: instructionEven = 32'h0;
	380: instructionEven = 32'h0;
	381: instructionEven = 32'h0;
	382: instructionEven = 32'h0;
	383: instructionEven = 32'h0;
	384: instructionEven = 32'h0;
	385: instructionEven = 32'h0;
	386: instructionEven = 32'h0;
	387: instructionEven = 32'h0;
	388: instructionEven = 32'h0;
	389: instructionEven = 32'h0;
	390: instructionEven = 32'h0;
	391: instructionEven = 32'h0;
	392: instructionEven = 32'h0;
	393: instructionEven = 32'h0;
	394: instructionEven = 32'h0;
	395: instructionEven = 32'h0;
	396: instructionEven = 32'h0;
	397: instructionEven = 32'h0;
	398: instructionEven = 32'h0;
	399: instructionEven = 32'h0;
	400: instructionEven = 32'h0;
	401: instructionEven = 32'h0;
	402: instructionEven = 32'h0;
	403: instructionEven = 32'h0;
	404: instructionEven = 32'h0;
	405: instructionEven = 32'h0;
	406: instructionEven = 32'h0;
	407: instructionEven = 32'h0;
	408: instructionEven = 32'h0;
	409: instructionEven = 32'h0;
	410: instructionEven = 32'h0;
	411: instructionEven = 32'h0;
	412: instructionEven = 32'h0;
	413: instructionEven = 32'h0;
	414: instructionEven = 32'h0;
	415: instructionEven = 32'h0;
	416: instructionEven = 32'h0;
	417: instructionEven = 32'h0;
	418: instructionEven = 32'h0;
	419: instructionEven = 32'h0;
	420: instructionEven = 32'h0;
	421: instructionEven = 32'h0;
	422: instructionEven = 32'h0;
	423: instructionEven = 32'h0;
	424: instructionEven = 32'h0;
	425: instructionEven = 32'h0;
	426: instructionEven = 32'h0;
	427: instructionEven = 32'h0;
	428: instructionEven = 32'h0;
	429: instructionEven = 32'h0;
	430: instructionEven = 32'h0;
	431: instructionEven = 32'h0;
	432: instructionEven = 32'h0;
	433: instructionEven = 32'h0;
	434: instructionEven = 32'h0;
	435: instructionEven = 32'h0;
	436: instructionEven = 32'h0;
	437: instructionEven = 32'h0;
	438: instructionEven = 32'h0;
	439: instructionEven = 32'h0;
	440: instructionEven = 32'h0;
	441: instructionEven = 32'h0;
	442: instructionEven = 32'h0;
	443: instructionEven = 32'h0;
	444: instructionEven = 32'h0;
	445: instructionEven = 32'h0;
	446: instructionEven = 32'h0;
	447: instructionEven = 32'h0;
	448: instructionEven = 32'h0;
	449: instructionEven = 32'h0;
	450: instructionEven = 32'h0;
	451: instructionEven = 32'h0;
	452: instructionEven = 32'h0;
	453: instructionEven = 32'h0;
	454: instructionEven = 32'h0;
	455: instructionEven = 32'h0;
	456: instructionEven = 32'h0;
	457: instructionEven = 32'h0;
	458: instructionEven = 32'h0;
	459: instructionEven = 32'h0;
	460: instructionEven = 32'h0;
	461: instructionEven = 32'h0;
	462: instructionEven = 32'h0;
	463: instructionEven = 32'h0;
	464: instructionEven = 32'h0;
	465: instructionEven = 32'h0;
	466: instructionEven = 32'h0;
	467: instructionEven = 32'h0;
	468: instructionEven = 32'h0;
	469: instructionEven = 32'h0;
	470: instructionEven = 32'h0;
	471: instructionEven = 32'h0;
	472: instructionEven = 32'h0;
	473: instructionEven = 32'h0;
	474: instructionEven = 32'h0;
	475: instructionEven = 32'h0;
	476: instructionEven = 32'h0;
	477: instructionEven = 32'h0;
	478: instructionEven = 32'h0;
	479: instructionEven = 32'h0;
	480: instructionEven = 32'h0;
	481: instructionEven = 32'h0;
	482: instructionEven = 32'h0;
	483: instructionEven = 32'h0;
	484: instructionEven = 32'h0;
	485: instructionEven = 32'h0;
	486: instructionEven = 32'h0;
	487: instructionEven = 32'h0;
	488: instructionEven = 32'h0;
	489: instructionEven = 32'h0;
	490: instructionEven = 32'h0;
	491: instructionEven = 32'h0;
	492: instructionEven = 32'h0;
	493: instructionEven = 32'h0;
	494: instructionEven = 32'h0;
	495: instructionEven = 32'h0;
	496: instructionEven = 32'h0;
	497: instructionEven = 32'h0;
	498: instructionEven = 32'h0;
	499: instructionEven = 32'h0;
	500: instructionEven = 32'h0;
	501: instructionEven = 32'h0;
	502: instructionEven = 32'h0;
	503: instructionEven = 32'h0;
	504: instructionEven = 32'h0;
	505: instructionEven = 32'h0;
	506: instructionEven = 32'h0;
	507: instructionEven = 32'h0;
	508: instructionEven = 32'h0;
	509: instructionEven = 32'h0;
	510: instructionEven = 32'h0;
	511: instructionEven = 32'h0;
	512: instructionEven = 32'h0;
	513: instructionEven = 32'h0;
	514: instructionEven = 32'h0;
	515: instructionEven = 32'h0;
	516: instructionEven = 32'h0;
	517: instructionEven = 32'h0;
	518: instructionEven = 32'h0;
	519: instructionEven = 32'h0;
	520: instructionEven = 32'h0;
	521: instructionEven = 32'h0;
	522: instructionEven = 32'h0;
	523: instructionEven = 32'h0;
	524: instructionEven = 32'h0;
	525: instructionEven = 32'h0;
	526: instructionEven = 32'h0;
	527: instructionEven = 32'h0;
	528: instructionEven = 32'h0;
	529: instructionEven = 32'h0;
	530: instructionEven = 32'h0;
	531: instructionEven = 32'h0;
	532: instructionEven = 32'h0;
	533: instructionEven = 32'h0;
	534: instructionEven = 32'h0;
	535: instructionEven = 32'h0;
	536: instructionEven = 32'h0;
	537: instructionEven = 32'h0;
	538: instructionEven = 32'h0;
	539: instructionEven = 32'h0;
	540: instructionEven = 32'h0;
	541: instructionEven = 32'h0;
	542: instructionEven = 32'h0;
	543: instructionEven = 32'h0;
	544: instructionEven = 32'h0;
	545: instructionEven = 32'h0;
	546: instructionEven = 32'h0;
	547: instructionEven = 32'h0;
	548: instructionEven = 32'h0;
	549: instructionEven = 32'h0;
	550: instructionEven = 32'h0;
	551: instructionEven = 32'h0;
	552: instructionEven = 32'h0;
	553: instructionEven = 32'h0;
	554: instructionEven = 32'h0;
	555: instructionEven = 32'h0;
	556: instructionEven = 32'h0;
	557: instructionEven = 32'h0;
	558: instructionEven = 32'h0;
	559: instructionEven = 32'h0;
	560: instructionEven = 32'h0;
	561: instructionEven = 32'h0;
	562: instructionEven = 32'h0;
	563: instructionEven = 32'h0;
	564: instructionEven = 32'h0;
	565: instructionEven = 32'h0;
	566: instructionEven = 32'h0;
	567: instructionEven = 32'h0;
	568: instructionEven = 32'h0;
	569: instructionEven = 32'h0;
	570: instructionEven = 32'h0;
	571: instructionEven = 32'h0;
	572: instructionEven = 32'h0;
	573: instructionEven = 32'h0;
	574: instructionEven = 32'h0;
	575: instructionEven = 32'h0;
	576: instructionEven = 32'h0;
	577: instructionEven = 32'h0;
	578: instructionEven = 32'h0;
	579: instructionEven = 32'h0;
	580: instructionEven = 32'h0;
	581: instructionEven = 32'h0;
	582: instructionEven = 32'h0;
	583: instructionEven = 32'h0;
	584: instructionEven = 32'h0;
	585: instructionEven = 32'h0;
	586: instructionEven = 32'h0;
	587: instructionEven = 32'h0;
	588: instructionEven = 32'h0;
	589: instructionEven = 32'h0;
	590: instructionEven = 32'h0;
	591: instructionEven = 32'h0;
	592: instructionEven = 32'h0;
	593: instructionEven = 32'h0;
	594: instructionEven = 32'h0;
	595: instructionEven = 32'h0;
	596: instructionEven = 32'h0;
	597: instructionEven = 32'h0;
	598: instructionEven = 32'h0;
	599: instructionEven = 32'h0;
	600: instructionEven = 32'h0;
	601: instructionEven = 32'h0;
	602: instructionEven = 32'h0;
	603: instructionEven = 32'h0;
	604: instructionEven = 32'h0;
	605: instructionEven = 32'h0;
	606: instructionEven = 32'h0;
	607: instructionEven = 32'h0;
	608: instructionEven = 32'h0;
	609: instructionEven = 32'h0;
	610: instructionEven = 32'h0;
	611: instructionEven = 32'h0;
	612: instructionEven = 32'h0;
	613: instructionEven = 32'h0;
	614: instructionEven = 32'h0;
	615: instructionEven = 32'h0;
	616: instructionEven = 32'h0;
	617: instructionEven = 32'h0;
	618: instructionEven = 32'h0;
	619: instructionEven = 32'h0;
	620: instructionEven = 32'h0;
	621: instructionEven = 32'h0;
	622: instructionEven = 32'h0;
	623: instructionEven = 32'h0;
	624: instructionEven = 32'h0;
	625: instructionEven = 32'h0;
	626: instructionEven = 32'h0;
	627: instructionEven = 32'h0;
	628: instructionEven = 32'h0;
	629: instructionEven = 32'h0;
	630: instructionEven = 32'h0;
	631: instructionEven = 32'h0;
	632: instructionEven = 32'h0;
	633: instructionEven = 32'h0;
	634: instructionEven = 32'h0;
	635: instructionEven = 32'h0;
	636: instructionEven = 32'h0;
	637: instructionEven = 32'h0;
	638: instructionEven = 32'h0;
	639: instructionEven = 32'h0;
	640: instructionEven = 32'h0;
	641: instructionEven = 32'h0;
	642: instructionEven = 32'h0;
	643: instructionEven = 32'h0;
	644: instructionEven = 32'h0;
	645: instructionEven = 32'h0;
	646: instructionEven = 32'h0;
	647: instructionEven = 32'h0;
	648: instructionEven = 32'h0;
	649: instructionEven = 32'h0;
	650: instructionEven = 32'h0;
	651: instructionEven = 32'h0;
	652: instructionEven = 32'h0;
	653: instructionEven = 32'h0;
	654: instructionEven = 32'h0;
	655: instructionEven = 32'h0;
	656: instructionEven = 32'h0;
	657: instructionEven = 32'h0;
	658: instructionEven = 32'h0;
	659: instructionEven = 32'h0;
	660: instructionEven = 32'h0;
	661: instructionEven = 32'h0;
	662: instructionEven = 32'h0;
	663: instructionEven = 32'h0;
	664: instructionEven = 32'h0;
	665: instructionEven = 32'h0;
	666: instructionEven = 32'h0;
	667: instructionEven = 32'h0;
	668: instructionEven = 32'h0;
	669: instructionEven = 32'h0;
	670: instructionEven = 32'h0;
	671: instructionEven = 32'h0;
	672: instructionEven = 32'h0;
	673: instructionEven = 32'h0;
	674: instructionEven = 32'h0;
	675: instructionEven = 32'h0;
	676: instructionEven = 32'h0;
	677: instructionEven = 32'h0;
	678: instructionEven = 32'h0;
	679: instructionEven = 32'h0;
	680: instructionEven = 32'h0;
	681: instructionEven = 32'h0;
	682: instructionEven = 32'h0;
	683: instructionEven = 32'h0;
	684: instructionEven = 32'h0;
	685: instructionEven = 32'h0;
	686: instructionEven = 32'h0;
	687: instructionEven = 32'h0;
	688: instructionEven = 32'h0;
	689: instructionEven = 32'h0;
	690: instructionEven = 32'h0;
	691: instructionEven = 32'h0;
	692: instructionEven = 32'h0;
	693: instructionEven = 32'h0;
	694: instructionEven = 32'h0;
	695: instructionEven = 32'h0;
	696: instructionEven = 32'h0;
	697: instructionEven = 32'h0;
	698: instructionEven = 32'h0;
	699: instructionEven = 32'h0;
	700: instructionEven = 32'h0;
	701: instructionEven = 32'h0;
	702: instructionEven = 32'h0;
	703: instructionEven = 32'h0;
	704: instructionEven = 32'h0;
	705: instructionEven = 32'h0;
	706: instructionEven = 32'h0;
	707: instructionEven = 32'h0;
	708: instructionEven = 32'h0;
	709: instructionEven = 32'h0;
	710: instructionEven = 32'h0;
	711: instructionEven = 32'h0;
	712: instructionEven = 32'h0;
	713: instructionEven = 32'h0;
	714: instructionEven = 32'h0;
	715: instructionEven = 32'h0;
	716: instructionEven = 32'h0;
	717: instructionEven = 32'h0;
	718: instructionEven = 32'h0;
	719: instructionEven = 32'h0;
	720: instructionEven = 32'h0;
	721: instructionEven = 32'h0;
	722: instructionEven = 32'h0;
	723: instructionEven = 32'h0;
	724: instructionEven = 32'h0;
	725: instructionEven = 32'h0;
	726: instructionEven = 32'h0;
	727: instructionEven = 32'h0;
	728: instructionEven = 32'h0;
	729: instructionEven = 32'h0;
	730: instructionEven = 32'h0;
	731: instructionEven = 32'h0;
	732: instructionEven = 32'h0;
	733: instructionEven = 32'h0;
	734: instructionEven = 32'h0;
	735: instructionEven = 32'h0;
	736: instructionEven = 32'h0;
	737: instructionEven = 32'h0;
	738: instructionEven = 32'h0;
	739: instructionEven = 32'h0;
	740: instructionEven = 32'h0;
	741: instructionEven = 32'h0;
	742: instructionEven = 32'h0;
	743: instructionEven = 32'h0;
	744: instructionEven = 32'h0;
	745: instructionEven = 32'h0;
	746: instructionEven = 32'h0;
	747: instructionEven = 32'h0;
	748: instructionEven = 32'h0;
	749: instructionEven = 32'h0;
	750: instructionEven = 32'h0;
	751: instructionEven = 32'h0;
	752: instructionEven = 32'h0;
	753: instructionEven = 32'h0;
	754: instructionEven = 32'h0;
	755: instructionEven = 32'h0;
	756: instructionEven = 32'h0;
	757: instructionEven = 32'h0;
	758: instructionEven = 32'h0;
	759: instructionEven = 32'h0;
	760: instructionEven = 32'h0;
	761: instructionEven = 32'h0;
	762: instructionEven = 32'h0;
	763: instructionEven = 32'h0;
	764: instructionEven = 32'h0;
	765: instructionEven = 32'h0;
	766: instructionEven = 32'h0;
	767: instructionEven = 32'h0;
	768: instructionEven = 32'h0;
	769: instructionEven = 32'h0;
	770: instructionEven = 32'h0;
	771: instructionEven = 32'h0;
	772: instructionEven = 32'h0;
	773: instructionEven = 32'h0;
	774: instructionEven = 32'h0;
	775: instructionEven = 32'h0;
	776: instructionEven = 32'h0;
	777: instructionEven = 32'h0;
	778: instructionEven = 32'h0;
	779: instructionEven = 32'h0;
	780: instructionEven = 32'h0;
	781: instructionEven = 32'h0;
	782: instructionEven = 32'h0;
	783: instructionEven = 32'h0;
	784: instructionEven = 32'h0;
	785: instructionEven = 32'h0;
	786: instructionEven = 32'h0;
	787: instructionEven = 32'h0;
	788: instructionEven = 32'h0;
	789: instructionEven = 32'h0;
	790: instructionEven = 32'h0;
	791: instructionEven = 32'h0;
	792: instructionEven = 32'h0;
	793: instructionEven = 32'h0;
	794: instructionEven = 32'h0;
	795: instructionEven = 32'h0;
	796: instructionEven = 32'h0;
	797: instructionEven = 32'h0;
	798: instructionEven = 32'h0;
	799: instructionEven = 32'h0;
	800: instructionEven = 32'h0;
	801: instructionEven = 32'h0;
	802: instructionEven = 32'h0;
	803: instructionEven = 32'h0;
	804: instructionEven = 32'h0;
	805: instructionEven = 32'h0;
	806: instructionEven = 32'h0;
	807: instructionEven = 32'h0;
	808: instructionEven = 32'h0;
	809: instructionEven = 32'h0;
	810: instructionEven = 32'h0;
	811: instructionEven = 32'h0;
	812: instructionEven = 32'h0;
	813: instructionEven = 32'h0;
	814: instructionEven = 32'h0;
	815: instructionEven = 32'h0;
	816: instructionEven = 32'h0;
	817: instructionEven = 32'h0;
	818: instructionEven = 32'h0;
	819: instructionEven = 32'h0;
	820: instructionEven = 32'h0;
	821: instructionEven = 32'h0;
	822: instructionEven = 32'h0;
	823: instructionEven = 32'h0;
	824: instructionEven = 32'h0;
	825: instructionEven = 32'h0;
	826: instructionEven = 32'h0;
	827: instructionEven = 32'h0;
	828: instructionEven = 32'h0;
	829: instructionEven = 32'h0;
	830: instructionEven = 32'h0;
	831: instructionEven = 32'h0;
	832: instructionEven = 32'h0;
	833: instructionEven = 32'h0;
	834: instructionEven = 32'h0;
	835: instructionEven = 32'h0;
	836: instructionEven = 32'h0;
	837: instructionEven = 32'h0;
	838: instructionEven = 32'h0;
	839: instructionEven = 32'h0;
	840: instructionEven = 32'h0;
	841: instructionEven = 32'h0;
	842: instructionEven = 32'h0;
	843: instructionEven = 32'h0;
	844: instructionEven = 32'h0;
	845: instructionEven = 32'h0;
	846: instructionEven = 32'h0;
	847: instructionEven = 32'h0;
	848: instructionEven = 32'h0;
	849: instructionEven = 32'h0;
	850: instructionEven = 32'h0;
	851: instructionEven = 32'h0;
	852: instructionEven = 32'h0;
	853: instructionEven = 32'h0;
	854: instructionEven = 32'h0;
	855: instructionEven = 32'h0;
	856: instructionEven = 32'h0;
	857: instructionEven = 32'h0;
	858: instructionEven = 32'h0;
	859: instructionEven = 32'h0;
	860: instructionEven = 32'h0;
	861: instructionEven = 32'h0;
	862: instructionEven = 32'h0;
	863: instructionEven = 32'h0;
	864: instructionEven = 32'h0;
	865: instructionEven = 32'h0;
	866: instructionEven = 32'h0;
	867: instructionEven = 32'h0;
	868: instructionEven = 32'h0;
	869: instructionEven = 32'h0;
	870: instructionEven = 32'h0;
	871: instructionEven = 32'h0;
	872: instructionEven = 32'h0;
	873: instructionEven = 32'h0;
	874: instructionEven = 32'h0;
	875: instructionEven = 32'h0;
	876: instructionEven = 32'h0;
	877: instructionEven = 32'h0;
	878: instructionEven = 32'h0;
	879: instructionEven = 32'h0;
	880: instructionEven = 32'h0;
	881: instructionEven = 32'h0;
	882: instructionEven = 32'h0;
	883: instructionEven = 32'h0;
	884: instructionEven = 32'h0;
	885: instructionEven = 32'h0;
	886: instructionEven = 32'h0;
	887: instructionEven = 32'h0;
	888: instructionEven = 32'h0;
	889: instructionEven = 32'h0;
	890: instructionEven = 32'h0;
	891: instructionEven = 32'h0;
	892: instructionEven = 32'h0;
	893: instructionEven = 32'h0;
	894: instructionEven = 32'h0;
	895: instructionEven = 32'h0;
	896: instructionEven = 32'h0;
	897: instructionEven = 32'h0;
	898: instructionEven = 32'h0;
	899: instructionEven = 32'h0;
	900: instructionEven = 32'h0;
	901: instructionEven = 32'h0;
	902: instructionEven = 32'h0;
	903: instructionEven = 32'h0;
	904: instructionEven = 32'h0;
	905: instructionEven = 32'h0;
	906: instructionEven = 32'h0;
	907: instructionEven = 32'h0;
	908: instructionEven = 32'h0;
	909: instructionEven = 32'h0;
	910: instructionEven = 32'h0;
	911: instructionEven = 32'h0;
	912: instructionEven = 32'h0;
	913: instructionEven = 32'h0;
	914: instructionEven = 32'h0;
	915: instructionEven = 32'h0;
	916: instructionEven = 32'h0;
	917: instructionEven = 32'h0;
	918: instructionEven = 32'h0;
	919: instructionEven = 32'h0;
	920: instructionEven = 32'h0;
	921: instructionEven = 32'h0;
	922: instructionEven = 32'h0;
	923: instructionEven = 32'h0;
	924: instructionEven = 32'h0;
	925: instructionEven = 32'h0;
	926: instructionEven = 32'h0;
	927: instructionEven = 32'h0;
	928: instructionEven = 32'h0;
	929: instructionEven = 32'h0;
	930: instructionEven = 32'h0;
	931: instructionEven = 32'h0;
	932: instructionEven = 32'h0;
	933: instructionEven = 32'h0;
	934: instructionEven = 32'h0;
	935: instructionEven = 32'h0;
	936: instructionEven = 32'h0;
	937: instructionEven = 32'h0;
	938: instructionEven = 32'h0;
	939: instructionEven = 32'h0;
	940: instructionEven = 32'h0;
	941: instructionEven = 32'h0;
	942: instructionEven = 32'h0;
	943: instructionEven = 32'h0;
	944: instructionEven = 32'h0;
	945: instructionEven = 32'h0;
	946: instructionEven = 32'h0;
	947: instructionEven = 32'h0;
	948: instructionEven = 32'h0;
	949: instructionEven = 32'h0;
	950: instructionEven = 32'h0;
	951: instructionEven = 32'h0;
	952: instructionEven = 32'h0;
	953: instructionEven = 32'h0;
	954: instructionEven = 32'h0;
	955: instructionEven = 32'h0;
	956: instructionEven = 32'h0;
	957: instructionEven = 32'h0;
	958: instructionEven = 32'h0;
	959: instructionEven = 32'h0;
	960: instructionEven = 32'h0;
	961: instructionEven = 32'h0;
	962: instructionEven = 32'h0;
	963: instructionEven = 32'h0;
	964: instructionEven = 32'h0;
	965: instructionEven = 32'h0;
	966: instructionEven = 32'h0;
	967: instructionEven = 32'h0;
	968: instructionEven = 32'h0;
	969: instructionEven = 32'h0;
	970: instructionEven = 32'h0;
	971: instructionEven = 32'h0;
	972: instructionEven = 32'h0;
	973: instructionEven = 32'h0;
	974: instructionEven = 32'h0;
	975: instructionEven = 32'h0;
	976: instructionEven = 32'h0;
	977: instructionEven = 32'h0;
	978: instructionEven = 32'h0;
	979: instructionEven = 32'h0;
	980: instructionEven = 32'h0;
	981: instructionEven = 32'h0;
	982: instructionEven = 32'h0;
	983: instructionEven = 32'h0;
	984: instructionEven = 32'h0;
	985: instructionEven = 32'h0;
	986: instructionEven = 32'h0;
	987: instructionEven = 32'h0;
	988: instructionEven = 32'h0;
	989: instructionEven = 32'h0;
	990: instructionEven = 32'h0;
	991: instructionEven = 32'h0;
	992: instructionEven = 32'h0;
	993: instructionEven = 32'h0;
	994: instructionEven = 32'h0;
	995: instructionEven = 32'h0;
	996: instructionEven = 32'h0;
	997: instructionEven = 32'h0;
	998: instructionEven = 32'h0;
	999: instructionEven = 32'h0;
	1000: instructionEven = 32'h0;
	1001: instructionEven = 32'h0;
	1002: instructionEven = 32'h0;
	1003: instructionEven = 32'h0;
	1004: instructionEven = 32'h0;
	1005: instructionEven = 32'h0;
	1006: instructionEven = 32'h0;
	1007: instructionEven = 32'h0;
	1008: instructionEven = 32'h0;
	1009: instructionEven = 32'h0;
	1010: instructionEven = 32'h0;
	1011: instructionEven = 32'h0;
	1012: instructionEven = 32'h0;
	1013: instructionEven = 32'h0;
	1014: instructionEven = 32'h0;
	1015: instructionEven = 32'h0;
	1016: instructionEven = 32'h0;
	1017: instructionEven = 32'h0;
	1018: instructionEven = 32'h0;
	1019: instructionEven = 32'h0;
	1020: instructionEven = 32'h0;
	1021: instructionEven = 32'h0;
	1022: instructionEven = 32'h0;
	1023: instructionEven = 32'h0;
	1024: instructionEven = 32'h0;
	1025: instructionEven = 32'h0;
	1026: instructionEven = 32'h0;
	1027: instructionEven = 32'h0;
	1028: instructionEven = 32'h0;
	1029: instructionEven = 32'h0;
	1030: instructionEven = 32'h0;
	1031: instructionEven = 32'h0;
	1032: instructionEven = 32'h0;
	1033: instructionEven = 32'h0;
	1034: instructionEven = 32'h0;
	1035: instructionEven = 32'h0;
	1036: instructionEven = 32'h0;
	1037: instructionEven = 32'h0;
	1038: instructionEven = 32'h0;
	1039: instructionEven = 32'h0;
	1040: instructionEven = 32'h0;
	1041: instructionEven = 32'h0;
	1042: instructionEven = 32'h0;
	1043: instructionEven = 32'h0;
	1044: instructionEven = 32'h0;
	1045: instructionEven = 32'h0;
	1046: instructionEven = 32'h0;
	1047: instructionEven = 32'h0;
	1048: instructionEven = 32'h0;
	1049: instructionEven = 32'h0;
	1050: instructionEven = 32'h0;
	1051: instructionEven = 32'h0;
	1052: instructionEven = 32'h0;
	1053: instructionEven = 32'h0;
	1054: instructionEven = 32'h0;
	1055: instructionEven = 32'h0;
	1056: instructionEven = 32'h0;
	1057: instructionEven = 32'h0;
	1058: instructionEven = 32'h0;
	1059: instructionEven = 32'h0;
	1060: instructionEven = 32'h0;
	1061: instructionEven = 32'h0;
	1062: instructionEven = 32'h0;
	1063: instructionEven = 32'h0;
	1064: instructionEven = 32'h0;
	1065: instructionEven = 32'h0;
	1066: instructionEven = 32'h0;
	1067: instructionEven = 32'h0;
	1068: instructionEven = 32'h0;
	1069: instructionEven = 32'h0;
	1070: instructionEven = 32'h0;
	1071: instructionEven = 32'h0;
	1072: instructionEven = 32'h0;
	1073: instructionEven = 32'h0;
	1074: instructionEven = 32'h0;
	1075: instructionEven = 32'h0;
	1076: instructionEven = 32'h0;
	1077: instructionEven = 32'h0;
	1078: instructionEven = 32'h0;
	1079: instructionEven = 32'h0;
	1080: instructionEven = 32'h0;
	1081: instructionEven = 32'h0;
	1082: instructionEven = 32'h0;
	1083: instructionEven = 32'h0;
	1084: instructionEven = 32'h0;
	1085: instructionEven = 32'h0;
	1086: instructionEven = 32'h0;
	1087: instructionEven = 32'h0;
	1088: instructionEven = 32'h0;
	1089: instructionEven = 32'h0;
	1090: instructionEven = 32'h0;
	1091: instructionEven = 32'h0;
	1092: instructionEven = 32'h0;
	1093: instructionEven = 32'h0;
	1094: instructionEven = 32'h0;
	1095: instructionEven = 32'h0;
	1096: instructionEven = 32'h0;
	1097: instructionEven = 32'h0;
	1098: instructionEven = 32'h0;
	1099: instructionEven = 32'h0;
	1100: instructionEven = 32'h0;
	1101: instructionEven = 32'h0;
	1102: instructionEven = 32'h0;
	1103: instructionEven = 32'h0;
	1104: instructionEven = 32'h0;
	1105: instructionEven = 32'h0;
	1106: instructionEven = 32'h0;
	1107: instructionEven = 32'h0;
	1108: instructionEven = 32'h0;
	1109: instructionEven = 32'h0;
	1110: instructionEven = 32'h0;
	1111: instructionEven = 32'h0;
	1112: instructionEven = 32'h0;
	1113: instructionEven = 32'h0;
	1114: instructionEven = 32'h0;
	1115: instructionEven = 32'h0;
	1116: instructionEven = 32'h0;
	1117: instructionEven = 32'h0;
	1118: instructionEven = 32'h0;
	1119: instructionEven = 32'h0;
	1120: instructionEven = 32'h0;
	1121: instructionEven = 32'h0;
	1122: instructionEven = 32'h0;
	1123: instructionEven = 32'h0;
	1124: instructionEven = 32'h0;
	1125: instructionEven = 32'h0;
	1126: instructionEven = 32'h0;
	1127: instructionEven = 32'h0;
	1128: instructionEven = 32'h0;
	1129: instructionEven = 32'h0;
	1130: instructionEven = 32'h0;
	1131: instructionEven = 32'h0;
	1132: instructionEven = 32'h0;
	1133: instructionEven = 32'h0;
	1134: instructionEven = 32'h0;
	1135: instructionEven = 32'h0;
	1136: instructionEven = 32'h0;
	1137: instructionEven = 32'h0;
	1138: instructionEven = 32'h0;
	1139: instructionEven = 32'h0;
	1140: instructionEven = 32'h0;
	1141: instructionEven = 32'h0;
	1142: instructionEven = 32'h0;
	1143: instructionEven = 32'h0;
	1144: instructionEven = 32'h0;
	1145: instructionEven = 32'h0;
	1146: instructionEven = 32'h0;
	1147: instructionEven = 32'h0;
	1148: instructionEven = 32'h0;
	1149: instructionEven = 32'h0;
	1150: instructionEven = 32'h0;
	1151: instructionEven = 32'h0;
	1152: instructionEven = 32'h0;
	1153: instructionEven = 32'h0;
	1154: instructionEven = 32'h0;
	1155: instructionEven = 32'h0;
	1156: instructionEven = 32'h0;
	1157: instructionEven = 32'h0;
	1158: instructionEven = 32'h0;
	1159: instructionEven = 32'h0;
	1160: instructionEven = 32'h0;
	1161: instructionEven = 32'h0;
	1162: instructionEven = 32'h0;
	1163: instructionEven = 32'h0;
	1164: instructionEven = 32'h0;
	1165: instructionEven = 32'h0;
	1166: instructionEven = 32'h0;
	1167: instructionEven = 32'h0;
	1168: instructionEven = 32'h0;
	1169: instructionEven = 32'h0;
	1170: instructionEven = 32'h0;
	1171: instructionEven = 32'h0;
	1172: instructionEven = 32'h0;
	1173: instructionEven = 32'h0;
	1174: instructionEven = 32'h0;
	1175: instructionEven = 32'h0;
	1176: instructionEven = 32'h0;
	1177: instructionEven = 32'h0;
	1178: instructionEven = 32'h0;
	1179: instructionEven = 32'h0;
	1180: instructionEven = 32'h0;
	1181: instructionEven = 32'h0;
	1182: instructionEven = 32'h0;
	1183: instructionEven = 32'h0;
	1184: instructionEven = 32'h0;
	1185: instructionEven = 32'h0;
	1186: instructionEven = 32'h0;
	1187: instructionEven = 32'h0;
	1188: instructionEven = 32'h0;
	1189: instructionEven = 32'h0;
	1190: instructionEven = 32'h0;
	1191: instructionEven = 32'h0;
	1192: instructionEven = 32'h0;
	1193: instructionEven = 32'h0;
	1194: instructionEven = 32'h0;
	1195: instructionEven = 32'h0;
	1196: instructionEven = 32'h0;
	1197: instructionEven = 32'h0;
	1198: instructionEven = 32'h0;
	1199: instructionEven = 32'h0;
	1200: instructionEven = 32'h0;
	1201: instructionEven = 32'h0;
	1202: instructionEven = 32'h0;
	1203: instructionEven = 32'h0;
	1204: instructionEven = 32'h0;
	1205: instructionEven = 32'h0;
	1206: instructionEven = 32'h0;
	1207: instructionEven = 32'h0;
	1208: instructionEven = 32'h0;
	1209: instructionEven = 32'h0;
	1210: instructionEven = 32'h0;
	1211: instructionEven = 32'h0;
	1212: instructionEven = 32'h0;
	1213: instructionEven = 32'h0;
	1214: instructionEven = 32'h0;
	1215: instructionEven = 32'h0;
	1216: instructionEven = 32'h0;
	1217: instructionEven = 32'h0;
	1218: instructionEven = 32'h0;
	1219: instructionEven = 32'h0;
	1220: instructionEven = 32'h0;
	1221: instructionEven = 32'h0;
	1222: instructionEven = 32'h0;
	1223: instructionEven = 32'h0;
	1224: instructionEven = 32'h0;
	1225: instructionEven = 32'h0;
	1226: instructionEven = 32'h0;
	1227: instructionEven = 32'h0;
	1228: instructionEven = 32'h0;
	1229: instructionEven = 32'h0;
	1230: instructionEven = 32'h0;
	1231: instructionEven = 32'h0;
	1232: instructionEven = 32'h0;
	1233: instructionEven = 32'h0;
	1234: instructionEven = 32'h0;
	1235: instructionEven = 32'h0;
	1236: instructionEven = 32'h0;
	1237: instructionEven = 32'h0;
	1238: instructionEven = 32'h0;
	1239: instructionEven = 32'h0;
	1240: instructionEven = 32'h0;
	1241: instructionEven = 32'h0;
	1242: instructionEven = 32'h0;
	1243: instructionEven = 32'h0;
	1244: instructionEven = 32'h0;
	1245: instructionEven = 32'h0;
	1246: instructionEven = 32'h0;
	1247: instructionEven = 32'h0;
	1248: instructionEven = 32'h0;
	1249: instructionEven = 32'h0;
	1250: instructionEven = 32'h0;
	1251: instructionEven = 32'h0;
	1252: instructionEven = 32'h0;
	1253: instructionEven = 32'h0;
	1254: instructionEven = 32'h0;
	1255: instructionEven = 32'h0;
	1256: instructionEven = 32'h0;
	1257: instructionEven = 32'h0;
	1258: instructionEven = 32'h0;
	1259: instructionEven = 32'h0;
	1260: instructionEven = 32'h0;
	1261: instructionEven = 32'h0;
	1262: instructionEven = 32'h0;
	1263: instructionEven = 32'h0;
	1264: instructionEven = 32'h0;
	1265: instructionEven = 32'h0;
	1266: instructionEven = 32'h0;
	1267: instructionEven = 32'h0;
	1268: instructionEven = 32'h0;
	1269: instructionEven = 32'h0;
	1270: instructionEven = 32'h0;
	1271: instructionEven = 32'h0;
	1272: instructionEven = 32'h0;
	1273: instructionEven = 32'h0;
	1274: instructionEven = 32'h0;
	1275: instructionEven = 32'h0;
	1276: instructionEven = 32'h0;
	1277: instructionEven = 32'h0;
	1278: instructionEven = 32'h0;
	1279: instructionEven = 32'h0;
	1280: instructionEven = 32'h0;
	1281: instructionEven = 32'h0;
	1282: instructionEven = 32'h0;
	1283: instructionEven = 32'h0;
	1284: instructionEven = 32'h0;
	1285: instructionEven = 32'h0;
	1286: instructionEven = 32'h0;
	1287: instructionEven = 32'h0;
	1288: instructionEven = 32'h0;
	1289: instructionEven = 32'h0;
	1290: instructionEven = 32'h0;
	1291: instructionEven = 32'h0;
	1292: instructionEven = 32'h0;
	1293: instructionEven = 32'h0;
	1294: instructionEven = 32'h0;
	1295: instructionEven = 32'h0;
	1296: instructionEven = 32'h0;
	1297: instructionEven = 32'h0;
	1298: instructionEven = 32'h0;
	1299: instructionEven = 32'h0;
	1300: instructionEven = 32'h0;
	1301: instructionEven = 32'h0;
	1302: instructionEven = 32'h0;
	1303: instructionEven = 32'h0;
	1304: instructionEven = 32'h0;
	1305: instructionEven = 32'h0;
	1306: instructionEven = 32'h0;
	1307: instructionEven = 32'h0;
	1308: instructionEven = 32'h0;
	1309: instructionEven = 32'h0;
	1310: instructionEven = 32'h0;
	1311: instructionEven = 32'h0;
	1312: instructionEven = 32'h0;
	1313: instructionEven = 32'h0;
	1314: instructionEven = 32'h0;
	1315: instructionEven = 32'h0;
	1316: instructionEven = 32'h0;
	1317: instructionEven = 32'h0;
	1318: instructionEven = 32'h0;
	1319: instructionEven = 32'h0;
	1320: instructionEven = 32'h0;
	1321: instructionEven = 32'h0;
	1322: instructionEven = 32'h0;
	1323: instructionEven = 32'h0;
	1324: instructionEven = 32'h0;
	1325: instructionEven = 32'h0;
	1326: instructionEven = 32'h0;
	1327: instructionEven = 32'h0;
	1328: instructionEven = 32'h0;
	1329: instructionEven = 32'h0;
	1330: instructionEven = 32'h0;
	1331: instructionEven = 32'h0;
	1332: instructionEven = 32'h0;
	1333: instructionEven = 32'h0;
	1334: instructionEven = 32'h0;
	1335: instructionEven = 32'h0;
	1336: instructionEven = 32'h0;
	1337: instructionEven = 32'h0;
	1338: instructionEven = 32'h0;
	1339: instructionEven = 32'h0;
	1340: instructionEven = 32'h0;
	1341: instructionEven = 32'h0;
	1342: instructionEven = 32'h0;
	1343: instructionEven = 32'h0;
	1344: instructionEven = 32'h0;
	1345: instructionEven = 32'h0;
	1346: instructionEven = 32'h0;
	1347: instructionEven = 32'h0;
	1348: instructionEven = 32'h0;
	1349: instructionEven = 32'h0;
	1350: instructionEven = 32'h0;
	1351: instructionEven = 32'h0;
	1352: instructionEven = 32'h0;
	1353: instructionEven = 32'h0;
	1354: instructionEven = 32'h0;
	1355: instructionEven = 32'h0;
	1356: instructionEven = 32'h0;
	1357: instructionEven = 32'h0;
	1358: instructionEven = 32'h0;
	1359: instructionEven = 32'h0;
	1360: instructionEven = 32'h0;
	1361: instructionEven = 32'h0;
	1362: instructionEven = 32'h0;
	1363: instructionEven = 32'h0;
	1364: instructionEven = 32'h0;
	1365: instructionEven = 32'h0;
	1366: instructionEven = 32'h0;
	1367: instructionEven = 32'h0;
	1368: instructionEven = 32'h0;
	1369: instructionEven = 32'h0;
	1370: instructionEven = 32'h0;
	1371: instructionEven = 32'h0;
	1372: instructionEven = 32'h0;
	1373: instructionEven = 32'h0;
	1374: instructionEven = 32'h0;
	1375: instructionEven = 32'h0;
	1376: instructionEven = 32'h0;
	1377: instructionEven = 32'h0;
	1378: instructionEven = 32'h0;
	1379: instructionEven = 32'h0;
	1380: instructionEven = 32'h0;
	1381: instructionEven = 32'h0;
	1382: instructionEven = 32'h0;
	1383: instructionEven = 32'h0;
	1384: instructionEven = 32'h0;
	1385: instructionEven = 32'h0;
	1386: instructionEven = 32'h0;
	1387: instructionEven = 32'h0;
	1388: instructionEven = 32'h0;
	1389: instructionEven = 32'h0;
	1390: instructionEven = 32'h0;
	1391: instructionEven = 32'h0;
	1392: instructionEven = 32'h0;
	1393: instructionEven = 32'h0;
	1394: instructionEven = 32'h0;
	1395: instructionEven = 32'h0;
	1396: instructionEven = 32'h0;
	1397: instructionEven = 32'h0;
	1398: instructionEven = 32'h0;
	1399: instructionEven = 32'h0;
	1400: instructionEven = 32'h0;
	1401: instructionEven = 32'h0;
	1402: instructionEven = 32'h0;
	1403: instructionEven = 32'h0;
	1404: instructionEven = 32'h0;
	1405: instructionEven = 32'h0;
	1406: instructionEven = 32'h0;
	1407: instructionEven = 32'h0;
	1408: instructionEven = 32'h0;
	1409: instructionEven = 32'h0;
	1410: instructionEven = 32'h0;
	1411: instructionEven = 32'h0;
	1412: instructionEven = 32'h0;
	1413: instructionEven = 32'h0;
	1414: instructionEven = 32'h0;
	1415: instructionEven = 32'h0;
	1416: instructionEven = 32'h0;
	1417: instructionEven = 32'h0;
	1418: instructionEven = 32'h0;
	1419: instructionEven = 32'h0;
	1420: instructionEven = 32'h0;
	1421: instructionEven = 32'h0;
	1422: instructionEven = 32'h0;
	1423: instructionEven = 32'h0;
	1424: instructionEven = 32'h0;
	1425: instructionEven = 32'h0;
	1426: instructionEven = 32'h0;
	1427: instructionEven = 32'h0;
	1428: instructionEven = 32'h0;
	1429: instructionEven = 32'h0;
	1430: instructionEven = 32'h0;
	1431: instructionEven = 32'h0;
	1432: instructionEven = 32'h0;
	1433: instructionEven = 32'h0;
	1434: instructionEven = 32'h0;
	1435: instructionEven = 32'h0;
	1436: instructionEven = 32'h0;
	1437: instructionEven = 32'h0;
	1438: instructionEven = 32'h0;
	1439: instructionEven = 32'h0;
	1440: instructionEven = 32'h0;
	1441: instructionEven = 32'h0;
	1442: instructionEven = 32'h0;
	1443: instructionEven = 32'h0;
	1444: instructionEven = 32'h0;
	1445: instructionEven = 32'h0;
	1446: instructionEven = 32'h0;
	1447: instructionEven = 32'h0;
	1448: instructionEven = 32'h0;
	1449: instructionEven = 32'h0;
	1450: instructionEven = 32'h0;
	1451: instructionEven = 32'h0;
	1452: instructionEven = 32'h0;
	1453: instructionEven = 32'h0;
	1454: instructionEven = 32'h0;
	1455: instructionEven = 32'h0;
	1456: instructionEven = 32'h0;
	1457: instructionEven = 32'h0;
	1458: instructionEven = 32'h0;
	1459: instructionEven = 32'h0;
	1460: instructionEven = 32'h0;
	1461: instructionEven = 32'h0;
	1462: instructionEven = 32'h0;
	1463: instructionEven = 32'h0;
	1464: instructionEven = 32'h0;
	1465: instructionEven = 32'h0;
	1466: instructionEven = 32'h0;
	1467: instructionEven = 32'h0;
	1468: instructionEven = 32'h0;
	1469: instructionEven = 32'h0;
	1470: instructionEven = 32'h0;
	1471: instructionEven = 32'h0;
	1472: instructionEven = 32'h0;
	1473: instructionEven = 32'h0;
	1474: instructionEven = 32'h0;
	1475: instructionEven = 32'h0;
	1476: instructionEven = 32'h0;
	1477: instructionEven = 32'h0;
	1478: instructionEven = 32'h0;
	1479: instructionEven = 32'h0;
	1480: instructionEven = 32'h0;
	1481: instructionEven = 32'h0;
	1482: instructionEven = 32'h0;
	1483: instructionEven = 32'h0;
	1484: instructionEven = 32'h0;
	1485: instructionEven = 32'h0;
	1486: instructionEven = 32'h0;
	1487: instructionEven = 32'h0;
	1488: instructionEven = 32'h0;
	1489: instructionEven = 32'h0;
	1490: instructionEven = 32'h0;
	1491: instructionEven = 32'h0;
	1492: instructionEven = 32'h0;
	1493: instructionEven = 32'h0;
	1494: instructionEven = 32'h0;
	1495: instructionEven = 32'h0;
	1496: instructionEven = 32'h0;
	1497: instructionEven = 32'h0;
	1498: instructionEven = 32'h0;
	1499: instructionEven = 32'h0;
	1500: instructionEven = 32'h0;
	1501: instructionEven = 32'h0;
	1502: instructionEven = 32'h0;
	1503: instructionEven = 32'h0;
	1504: instructionEven = 32'h0;
	1505: instructionEven = 32'h0;
	1506: instructionEven = 32'h0;
	1507: instructionEven = 32'h0;
	1508: instructionEven = 32'h0;
	1509: instructionEven = 32'h0;
	1510: instructionEven = 32'h0;
	1511: instructionEven = 32'h0;
	1512: instructionEven = 32'h0;
	1513: instructionEven = 32'h0;
	1514: instructionEven = 32'h0;
	1515: instructionEven = 32'h0;
	1516: instructionEven = 32'h0;
	1517: instructionEven = 32'h0;
	1518: instructionEven = 32'h0;
	1519: instructionEven = 32'h0;
	1520: instructionEven = 32'h0;
	1521: instructionEven = 32'h0;
	1522: instructionEven = 32'h0;
	1523: instructionEven = 32'h0;
	1524: instructionEven = 32'h0;
	1525: instructionEven = 32'h0;
	1526: instructionEven = 32'h0;
	1527: instructionEven = 32'h0;
	1528: instructionEven = 32'h0;
	1529: instructionEven = 32'h0;
	1530: instructionEven = 32'h0;
	1531: instructionEven = 32'h0;
	1532: instructionEven = 32'h0;
	1533: instructionEven = 32'h0;
	1534: instructionEven = 32'h0;
	1535: instructionEven = 32'h0;
	1536: instructionEven = 32'h0;
	1537: instructionEven = 32'h0;
	1538: instructionEven = 32'h0;
	1539: instructionEven = 32'h0;
	1540: instructionEven = 32'h0;
	1541: instructionEven = 32'h0;
	1542: instructionEven = 32'h0;
	1543: instructionEven = 32'h0;
	1544: instructionEven = 32'h0;
	1545: instructionEven = 32'h0;
	1546: instructionEven = 32'h0;
	1547: instructionEven = 32'h0;
	1548: instructionEven = 32'h0;
	1549: instructionEven = 32'h0;
	1550: instructionEven = 32'h0;
	1551: instructionEven = 32'h0;
	1552: instructionEven = 32'h0;
	1553: instructionEven = 32'h0;
	1554: instructionEven = 32'h0;
	1555: instructionEven = 32'h0;
	1556: instructionEven = 32'h0;
	1557: instructionEven = 32'h0;
	1558: instructionEven = 32'h0;
	1559: instructionEven = 32'h0;
	1560: instructionEven = 32'h0;
	1561: instructionEven = 32'h0;
	1562: instructionEven = 32'h0;
	1563: instructionEven = 32'h0;
	1564: instructionEven = 32'h0;
	1565: instructionEven = 32'h0;
	1566: instructionEven = 32'h0;
	1567: instructionEven = 32'h0;
	1568: instructionEven = 32'h0;
	1569: instructionEven = 32'h0;
	1570: instructionEven = 32'h0;
	1571: instructionEven = 32'h0;
	1572: instructionEven = 32'h0;
	1573: instructionEven = 32'h0;
	1574: instructionEven = 32'h0;
	1575: instructionEven = 32'h0;
	1576: instructionEven = 32'h0;
	1577: instructionEven = 32'h0;
	1578: instructionEven = 32'h0;
	1579: instructionEven = 32'h0;
	1580: instructionEven = 32'h0;
	1581: instructionEven = 32'h0;
	1582: instructionEven = 32'h0;
	1583: instructionEven = 32'h0;
	1584: instructionEven = 32'h0;
	1585: instructionEven = 32'h0;
	1586: instructionEven = 32'h0;
	1587: instructionEven = 32'h0;
	1588: instructionEven = 32'h0;
	1589: instructionEven = 32'h0;
	1590: instructionEven = 32'h0;
	1591: instructionEven = 32'h0;
	1592: instructionEven = 32'h0;
	1593: instructionEven = 32'h0;
	1594: instructionEven = 32'h0;
	1595: instructionEven = 32'h0;
	1596: instructionEven = 32'h0;
	1597: instructionEven = 32'h0;
	1598: instructionEven = 32'h0;
	1599: instructionEven = 32'h0;
	1600: instructionEven = 32'h0;
	1601: instructionEven = 32'h0;
	1602: instructionEven = 32'h0;
	1603: instructionEven = 32'h0;
	1604: instructionEven = 32'h0;
	1605: instructionEven = 32'h0;
	1606: instructionEven = 32'h0;
	1607: instructionEven = 32'h0;
	1608: instructionEven = 32'h0;
	1609: instructionEven = 32'h0;
	1610: instructionEven = 32'h0;
	1611: instructionEven = 32'h0;
	1612: instructionEven = 32'h0;
	1613: instructionEven = 32'h0;
	1614: instructionEven = 32'h0;
	1615: instructionEven = 32'h0;
	1616: instructionEven = 32'h0;
	1617: instructionEven = 32'h0;
	1618: instructionEven = 32'h0;
	1619: instructionEven = 32'h0;
	1620: instructionEven = 32'h0;
	1621: instructionEven = 32'h0;
	1622: instructionEven = 32'h0;
	1623: instructionEven = 32'h0;
	1624: instructionEven = 32'h0;
	1625: instructionEven = 32'h0;
	1626: instructionEven = 32'h0;
	1627: instructionEven = 32'h0;
	1628: instructionEven = 32'h0;
	1629: instructionEven = 32'h0;
	1630: instructionEven = 32'h0;
	1631: instructionEven = 32'h0;
	1632: instructionEven = 32'h0;
	1633: instructionEven = 32'h0;
	1634: instructionEven = 32'h0;
	1635: instructionEven = 32'h0;
	1636: instructionEven = 32'h0;
	1637: instructionEven = 32'h0;
	1638: instructionEven = 32'h0;
	1639: instructionEven = 32'h0;
	1640: instructionEven = 32'h0;
	1641: instructionEven = 32'h0;
	1642: instructionEven = 32'h0;
	1643: instructionEven = 32'h0;
	1644: instructionEven = 32'h0;
	1645: instructionEven = 32'h0;
	1646: instructionEven = 32'h0;
	1647: instructionEven = 32'h0;
	1648: instructionEven = 32'h0;
	1649: instructionEven = 32'h0;
	1650: instructionEven = 32'h0;
	1651: instructionEven = 32'h0;
	1652: instructionEven = 32'h0;
	1653: instructionEven = 32'h0;
	1654: instructionEven = 32'h0;
	1655: instructionEven = 32'h0;
	1656: instructionEven = 32'h0;
	1657: instructionEven = 32'h0;
	1658: instructionEven = 32'h0;
	1659: instructionEven = 32'h0;
	1660: instructionEven = 32'h0;
	1661: instructionEven = 32'h0;
	1662: instructionEven = 32'h0;
	1663: instructionEven = 32'h0;
	1664: instructionEven = 32'h0;
	1665: instructionEven = 32'h0;
	1666: instructionEven = 32'h0;
	1667: instructionEven = 32'h0;
	1668: instructionEven = 32'h0;
	1669: instructionEven = 32'h0;
	1670: instructionEven = 32'h0;
	1671: instructionEven = 32'h0;
	1672: instructionEven = 32'h0;
	1673: instructionEven = 32'h0;
	1674: instructionEven = 32'h0;
	1675: instructionEven = 32'h0;
	1676: instructionEven = 32'h0;
	1677: instructionEven = 32'h0;
	1678: instructionEven = 32'h0;
	1679: instructionEven = 32'h0;
	1680: instructionEven = 32'h0;
	1681: instructionEven = 32'h0;
	1682: instructionEven = 32'h0;
	1683: instructionEven = 32'h0;
	1684: instructionEven = 32'h0;
	1685: instructionEven = 32'h0;
	1686: instructionEven = 32'h0;
	1687: instructionEven = 32'h0;
	1688: instructionEven = 32'h0;
	1689: instructionEven = 32'h0;
	1690: instructionEven = 32'h0;
	1691: instructionEven = 32'h0;
	1692: instructionEven = 32'h0;
	1693: instructionEven = 32'h0;
	1694: instructionEven = 32'h0;
	1695: instructionEven = 32'h0;
	1696: instructionEven = 32'h0;
	1697: instructionEven = 32'h0;
	1698: instructionEven = 32'h0;
	1699: instructionEven = 32'h0;
	1700: instructionEven = 32'h0;
	1701: instructionEven = 32'h0;
	1702: instructionEven = 32'h0;
	1703: instructionEven = 32'h0;
	1704: instructionEven = 32'h0;
	1705: instructionEven = 32'h0;
	1706: instructionEven = 32'h0;
	1707: instructionEven = 32'h0;
	1708: instructionEven = 32'h0;
	1709: instructionEven = 32'h0;
	1710: instructionEven = 32'h0;
	1711: instructionEven = 32'h0;
	1712: instructionEven = 32'h0;
	1713: instructionEven = 32'h0;
	1714: instructionEven = 32'h0;
	1715: instructionEven = 32'h0;
	1716: instructionEven = 32'h0;
	1717: instructionEven = 32'h0;
	1718: instructionEven = 32'h0;
	1719: instructionEven = 32'h0;
	1720: instructionEven = 32'h0;
	1721: instructionEven = 32'h0;
	1722: instructionEven = 32'h0;
	1723: instructionEven = 32'h0;
	1724: instructionEven = 32'h0;
	1725: instructionEven = 32'h0;
	1726: instructionEven = 32'h0;
	1727: instructionEven = 32'h0;
	1728: instructionEven = 32'h0;
	1729: instructionEven = 32'h0;
	1730: instructionEven = 32'h0;
	1731: instructionEven = 32'h0;
	1732: instructionEven = 32'h0;
	1733: instructionEven = 32'h0;
	1734: instructionEven = 32'h0;
	1735: instructionEven = 32'h0;
	1736: instructionEven = 32'h0;
	1737: instructionEven = 32'h0;
	1738: instructionEven = 32'h0;
	1739: instructionEven = 32'h0;
	1740: instructionEven = 32'h0;
	1741: instructionEven = 32'h0;
	1742: instructionEven = 32'h0;
	1743: instructionEven = 32'h0;
	1744: instructionEven = 32'h0;
	1745: instructionEven = 32'h0;
	1746: instructionEven = 32'h0;
	1747: instructionEven = 32'h0;
	1748: instructionEven = 32'h0;
	1749: instructionEven = 32'h0;
	1750: instructionEven = 32'h0;
	1751: instructionEven = 32'h0;
	1752: instructionEven = 32'h0;
	1753: instructionEven = 32'h0;
	1754: instructionEven = 32'h0;
	1755: instructionEven = 32'h0;
	1756: instructionEven = 32'h0;
	1757: instructionEven = 32'h0;
	1758: instructionEven = 32'h0;
	1759: instructionEven = 32'h0;
	1760: instructionEven = 32'h0;
	1761: instructionEven = 32'h0;
	1762: instructionEven = 32'h0;
	1763: instructionEven = 32'h0;
	1764: instructionEven = 32'h0;
	1765: instructionEven = 32'h0;
	1766: instructionEven = 32'h0;
	1767: instructionEven = 32'h0;
	1768: instructionEven = 32'h0;
	1769: instructionEven = 32'h0;
	1770: instructionEven = 32'h0;
	1771: instructionEven = 32'h0;
	1772: instructionEven = 32'h0;
	1773: instructionEven = 32'h0;
	1774: instructionEven = 32'h0;
	1775: instructionEven = 32'h0;
	1776: instructionEven = 32'h0;
	1777: instructionEven = 32'h0;
	1778: instructionEven = 32'h0;
	1779: instructionEven = 32'h0;
	1780: instructionEven = 32'h0;
	1781: instructionEven = 32'h0;
	1782: instructionEven = 32'h0;
	1783: instructionEven = 32'h0;
	1784: instructionEven = 32'h0;
	1785: instructionEven = 32'h0;
	1786: instructionEven = 32'h0;
	1787: instructionEven = 32'h0;
	1788: instructionEven = 32'h0;
	1789: instructionEven = 32'h0;
	1790: instructionEven = 32'h0;
	1791: instructionEven = 32'h0;
	1792: instructionEven = 32'h0;
	1793: instructionEven = 32'h0;
	1794: instructionEven = 32'h0;
	1795: instructionEven = 32'h0;
	1796: instructionEven = 32'h0;
	1797: instructionEven = 32'h0;
	1798: instructionEven = 32'h0;
	1799: instructionEven = 32'h0;
	1800: instructionEven = 32'h0;
	1801: instructionEven = 32'h0;
	1802: instructionEven = 32'h0;
	1803: instructionEven = 32'h0;
	1804: instructionEven = 32'h0;
	1805: instructionEven = 32'h0;
	1806: instructionEven = 32'h0;
	1807: instructionEven = 32'h0;
	1808: instructionEven = 32'h0;
	1809: instructionEven = 32'h0;
	1810: instructionEven = 32'h0;
	1811: instructionEven = 32'h0;
	1812: instructionEven = 32'h0;
	1813: instructionEven = 32'h0;
	1814: instructionEven = 32'h0;
	1815: instructionEven = 32'h0;
	1816: instructionEven = 32'h0;
	1817: instructionEven = 32'h0;
	1818: instructionEven = 32'h0;
	1819: instructionEven = 32'h0;
	1820: instructionEven = 32'h0;
	1821: instructionEven = 32'h0;
	1822: instructionEven = 32'h0;
	1823: instructionEven = 32'h0;
	1824: instructionEven = 32'h0;
	1825: instructionEven = 32'h0;
	1826: instructionEven = 32'h0;
	1827: instructionEven = 32'h0;
	1828: instructionEven = 32'h0;
	1829: instructionEven = 32'h0;
	1830: instructionEven = 32'h0;
	1831: instructionEven = 32'h0;
	1832: instructionEven = 32'h0;
	1833: instructionEven = 32'h0;
	1834: instructionEven = 32'h0;
	1835: instructionEven = 32'h0;
	1836: instructionEven = 32'h0;
	1837: instructionEven = 32'h0;
	1838: instructionEven = 32'h0;
	1839: instructionEven = 32'h0;
	1840: instructionEven = 32'h0;
	1841: instructionEven = 32'h0;
	1842: instructionEven = 32'h0;
	1843: instructionEven = 32'h0;
	1844: instructionEven = 32'h0;
	1845: instructionEven = 32'h0;
	1846: instructionEven = 32'h0;
	1847: instructionEven = 32'h0;
	1848: instructionEven = 32'h0;
	1849: instructionEven = 32'h0;
	1850: instructionEven = 32'h0;
	1851: instructionEven = 32'h0;
	1852: instructionEven = 32'h0;
	1853: instructionEven = 32'h0;
	1854: instructionEven = 32'h0;
	1855: instructionEven = 32'h0;
	1856: instructionEven = 32'h0;
	1857: instructionEven = 32'h0;
	1858: instructionEven = 32'h0;
	1859: instructionEven = 32'h0;
	1860: instructionEven = 32'h0;
	1861: instructionEven = 32'h0;
	1862: instructionEven = 32'h0;
	1863: instructionEven = 32'h0;
	1864: instructionEven = 32'h0;
	1865: instructionEven = 32'h0;
	1866: instructionEven = 32'h0;
	1867: instructionEven = 32'h0;
	1868: instructionEven = 32'h0;
	1869: instructionEven = 32'h0;
	1870: instructionEven = 32'h0;
	1871: instructionEven = 32'h0;
	1872: instructionEven = 32'h0;
	1873: instructionEven = 32'h0;
	1874: instructionEven = 32'h0;
	1875: instructionEven = 32'h0;
	1876: instructionEven = 32'h0;
	1877: instructionEven = 32'h0;
	1878: instructionEven = 32'h0;
	1879: instructionEven = 32'h0;
	1880: instructionEven = 32'h0;
	1881: instructionEven = 32'h0;
	1882: instructionEven = 32'h0;
	1883: instructionEven = 32'h0;
	1884: instructionEven = 32'h0;
	1885: instructionEven = 32'h0;
	1886: instructionEven = 32'h0;
	1887: instructionEven = 32'h0;
	1888: instructionEven = 32'h0;
	1889: instructionEven = 32'h0;
	1890: instructionEven = 32'h0;
	1891: instructionEven = 32'h0;
	1892: instructionEven = 32'h0;
	1893: instructionEven = 32'h0;
	1894: instructionEven = 32'h0;
	1895: instructionEven = 32'h0;
	1896: instructionEven = 32'h0;
	1897: instructionEven = 32'h0;
	1898: instructionEven = 32'h0;
	1899: instructionEven = 32'h0;
	1900: instructionEven = 32'h0;
	1901: instructionEven = 32'h0;
	1902: instructionEven = 32'h0;
	1903: instructionEven = 32'h0;
	1904: instructionEven = 32'h0;
	1905: instructionEven = 32'h0;
	1906: instructionEven = 32'h0;
	1907: instructionEven = 32'h0;
	1908: instructionEven = 32'h0;
	1909: instructionEven = 32'h0;
	1910: instructionEven = 32'h0;
	1911: instructionEven = 32'h0;
	1912: instructionEven = 32'h0;
	1913: instructionEven = 32'h0;
	1914: instructionEven = 32'h0;
	1915: instructionEven = 32'h0;
	1916: instructionEven = 32'h0;
	1917: instructionEven = 32'h0;
	1918: instructionEven = 32'h0;
	1919: instructionEven = 32'h0;
	1920: instructionEven = 32'h0;
	1921: instructionEven = 32'h0;
	1922: instructionEven = 32'h0;
	1923: instructionEven = 32'h0;
	1924: instructionEven = 32'h0;
	1925: instructionEven = 32'h0;
	1926: instructionEven = 32'h0;
	1927: instructionEven = 32'h0;
	1928: instructionEven = 32'h0;
	1929: instructionEven = 32'h0;
	1930: instructionEven = 32'h0;
	1931: instructionEven = 32'h0;
	1932: instructionEven = 32'h0;
	1933: instructionEven = 32'h0;
	1934: instructionEven = 32'h0;
	1935: instructionEven = 32'h0;
	1936: instructionEven = 32'h0;
	1937: instructionEven = 32'h0;
	1938: instructionEven = 32'h0;
	1939: instructionEven = 32'h0;
	1940: instructionEven = 32'h0;
	1941: instructionEven = 32'h0;
	1942: instructionEven = 32'h0;
	1943: instructionEven = 32'h0;
	1944: instructionEven = 32'h0;
	1945: instructionEven = 32'h0;
	1946: instructionEven = 32'h0;
	1947: instructionEven = 32'h0;
	1948: instructionEven = 32'h0;
	1949: instructionEven = 32'h0;
	1950: instructionEven = 32'h0;
	1951: instructionEven = 32'h0;
	1952: instructionEven = 32'h0;
	1953: instructionEven = 32'h0;
	1954: instructionEven = 32'h0;
	1955: instructionEven = 32'h0;
	1956: instructionEven = 32'h0;
	1957: instructionEven = 32'h0;
	1958: instructionEven = 32'h0;
	1959: instructionEven = 32'h0;
	1960: instructionEven = 32'h0;
	1961: instructionEven = 32'h0;
	1962: instructionEven = 32'h0;
	1963: instructionEven = 32'h0;
	1964: instructionEven = 32'h0;
	1965: instructionEven = 32'h0;
	1966: instructionEven = 32'h0;
	1967: instructionEven = 32'h0;
	1968: instructionEven = 32'h0;
	1969: instructionEven = 32'h0;
	1970: instructionEven = 32'h0;
	1971: instructionEven = 32'h0;
	1972: instructionEven = 32'h0;
	1973: instructionEven = 32'h0;
	1974: instructionEven = 32'h0;
	1975: instructionEven = 32'h0;
	1976: instructionEven = 32'h0;
	1977: instructionEven = 32'h0;
	1978: instructionEven = 32'h0;
	1979: instructionEven = 32'h0;
	1980: instructionEven = 32'h0;
	1981: instructionEven = 32'h0;
	1982: instructionEven = 32'h0;
	1983: instructionEven = 32'h0;
	1984: instructionEven = 32'h0;
	1985: instructionEven = 32'h0;
	1986: instructionEven = 32'h0;
	1987: instructionEven = 32'h0;
	1988: instructionEven = 32'h0;
	1989: instructionEven = 32'h0;
	1990: instructionEven = 32'h0;
	1991: instructionEven = 32'h0;
	1992: instructionEven = 32'h0;
	1993: instructionEven = 32'h0;
	1994: instructionEven = 32'h0;
	1995: instructionEven = 32'h0;
	1996: instructionEven = 32'h0;
	1997: instructionEven = 32'h0;
	1998: instructionEven = 32'h0;
	1999: instructionEven = 32'h0;
	2000: instructionEven = 32'h0;
	2001: instructionEven = 32'h0;
	2002: instructionEven = 32'h0;
	2003: instructionEven = 32'h0;
	2004: instructionEven = 32'h0;
	2005: instructionEven = 32'h0;
	2006: instructionEven = 32'h0;
	2007: instructionEven = 32'h0;
	2008: instructionEven = 32'h0;
	2009: instructionEven = 32'h0;
	2010: instructionEven = 32'h0;
	2011: instructionEven = 32'h0;
	2012: instructionEven = 32'h0;
	2013: instructionEven = 32'h0;
	2014: instructionEven = 32'h0;
	2015: instructionEven = 32'h0;
	2016: instructionEven = 32'h0;
	2017: instructionEven = 32'h0;
	2018: instructionEven = 32'h0;
	2019: instructionEven = 32'h0;
	2020: instructionEven = 32'h0;
	2021: instructionEven = 32'h0;
	2022: instructionEven = 32'h0;
	2023: instructionEven = 32'h0;
	2024: instructionEven = 32'h0;
	2025: instructionEven = 32'h0;
	2026: instructionEven = 32'h0;
	2027: instructionEven = 32'h0;
	2028: instructionEven = 32'h0;
	2029: instructionEven = 32'h0;
	2030: instructionEven = 32'h0;
	2031: instructionEven = 32'h0;
	2032: instructionEven = 32'h0;
	2033: instructionEven = 32'h0;
	2034: instructionEven = 32'h0;
	2035: instructionEven = 32'h0;
	2036: instructionEven = 32'h0;
	2037: instructionEven = 32'h0;
	2038: instructionEven = 32'h0;
	2039: instructionEven = 32'h0;
	2040: instructionEven = 32'h0;
	2041: instructionEven = 32'h0;
	2042: instructionEven = 32'h0;
	2043: instructionEven = 32'h0;
	2044: instructionEven = 32'h0;
	2045: instructionEven = 32'h0;
	2046: instructionEven = 32'h0;
	2047: instructionEven = 32'h0;

    default: begin
        instructionEven = 32'bx;
        `ifndef SYNTHESIS
            // synthesis translate_off
            instructionEven = {1{$random}};
            // synthesis translate_on
        `endif
    end
endcase
        
always @(*) case (addressOdd)
	0: instructionOdd = 32'h87c20000;
	1: instructionOdd = 32'h87c40000;
	2: instructionOdd = 32'h3e1000;
	3: instructionOdd = 32'h2402026;
	4: instructionOdd = 32'hf0010000;
	5: instructionOdd = 32'h400000;
	6: instructionOdd = 32'hcfc40000;
	7: instructionOdd = 32'hcfc20000;
	8: instructionOdd = 32'h4ac22085;
	9: instructionOdd = 32'h400000;
	10: instructionOdd = 32'h4800000;
	11: instructionOdd = 32'h7ff024;
	12: instructionOdd = 32'h2c5f482;
	13: instructionOdd = 32'h2520037;
	14: instructionOdd = 32'h2520030;
	15: instructionOdd = 32'h2c5fa83;
	16: instructionOdd = 32'h2c5fb85;
	17: instructionOdd = 32'h2c5fc87;
	18: instructionOdd = 32'hf0020000;
	19: instructionOdd = 32'h4403e8;
	20: instructionOdd = 32'h87c40000;
	21: instructionOdd = 32'h2842083;
	22: instructionOdd = 32'h2041100;
	23: instructionOdd = 32'hcbffffa;
	24: instructionOdd = 32'h2c60004;
	25: instructionOdd = 32'hf0000000;
	26: instructionOdd = 32'h400000;
	27: instructionOdd = 32'h4c800023;
	28: instructionOdd = 32'hf0000000;
	29: instructionOdd = 32'h400000;
	30: instructionOdd = 32'h2c62009;
	31: instructionOdd = 32'h460001;
	32: instructionOdd = 32'h2c62188;
	33: instructionOdd = 32'h400000;
	34: instructionOdd = 32'h2c62007;
	35: instructionOdd = 32'h400000;
	36: instructionOdd = 32'h2c61006;
	37: instructionOdd = 32'h87c20000;
	38: instructionOdd = 32'h2821080;
	39: instructionOdd = 32'hc21004;
	40: instructionOdd = 32'h2820185;
	41: instructionOdd = 32'h20210e1;
	42: instructionOdd = 32'h2820185;
	43: instructionOdd = 32'h2021161;
	44: instructionOdd = 32'h480001d;
	45: instructionOdd = 32'hf0000000;
	46: instructionOdd = 32'h400000;
	47: instructionOdd = 32'hcc00010;
	48: instructionOdd = 32'h40000;
	49: instructionOdd = 32'h2c61009;
	50: instructionOdd = 32'h2c61188;
	51: instructionOdd = 32'h2c61006;
	52: instructionOdd = 32'h87c60000;
	53: instructionOdd = 32'h2863082;
	54: instructionOdd = 32'h20221b4;
	55: instructionOdd = 32'h421001;
	56: instructionOdd = 32'hcfffffe;
	57: instructionOdd = 32'h2c60105;
	58: instructionOdd = 32'h2c60084;
	59: instructionOdd = 32'hf0000000;
	60: instructionOdd = 32'h400000;
	61: instructionOdd = 32'h20000;
	62: instructionOdd = 32'h87c4100d;
	63: instructionOdd = 32'h2862180;
	64: instructionOdd = 32'h2c22180;
	65: instructionOdd = 32'hf0000000;
	66: instructionOdd = 32'h21001;
	67: instructionOdd = 32'h2021134;
	68: instructionOdd = 32'h87c20000;
	69: instructionOdd = 32'h2821080;
	70: instructionOdd = 32'h2021031;
	71: instructionOdd = 32'h87c20000;
	72: instructionOdd = 32'h2821080;
	73: instructionOdd = 32'h4c00016;
	74: instructionOdd = 32'h2c61109;
	75: instructionOdd = 32'h2c60085;
	76: instructionOdd = 32'hf0000000;
	77: instructionOdd = 32'h20001;
	78: instructionOdd = 32'hc80000c;
	79: instructionOdd = 32'h2842189;
	80: instructionOdd = 32'h2022161;
	81: instructionOdd = 32'h87c40000;
	82: instructionOdd = 32'h2842082;
	83: instructionOdd = 32'h2021134;
	84: instructionOdd = 32'h2840184;
	85: instructionOdd = 32'h2022060;
	86: instructionOdd = 32'h87c20000;
	87: instructionOdd = 32'h2821085;
	88: instructionOdd = 32'h20220b2;
	89: instructionOdd = 32'hf0010000;
	90: instructionOdd = 32'h80000000;
	91: instructionOdd = 32'h400000;
	92: instructionOdd = 32'h2820184;
	93: instructionOdd = 32'h6001004;
	94: instructionOdd = 32'hf0010000;
	95: instructionOdd = 32'h400000;
	96: instructionOdd = 32'hcfc60000;
	97: instructionOdd = 32'hcfc40000;
	98: instructionOdd = 32'h4ac23105;
	99: instructionOdd = 32'h400000;
	100: instructionOdd = 32'hf0000000;
	101: instructionOdd = 32'h400000;
	102: instructionOdd = 32'h2c62088;
	103: instructionOdd = 32'h87c40000;
	104: instructionOdd = 32'h2842080;
	105: instructionOdd = 32'h2022031;
	106: instructionOdd = 32'h40004;
	107: instructionOdd = 32'hf0000000;
	108: instructionOdd = 32'h400000;
	109: instructionOdd = 32'h2c61109;
	110: instructionOdd = 32'h400000;
	111: instructionOdd = 32'hcbffff7;
	112: instructionOdd = 32'hf0000000;
	113: instructionOdd = 32'h4c00048;
	114: instructionOdd = 32'h2c61009;
	115: instructionOdd = 32'hf0000000;
	116: instructionOdd = 32'h40001;
	117: instructionOdd = 32'hc800011;
	118: instructionOdd = 32'h2863189;
	119: instructionOdd = 32'h2023060;
	120: instructionOdd = 32'hc62004;
	121: instructionOdd = 32'h400000;
	122: instructionOdd = 32'hcbffffc;
	123: instructionOdd = 32'hf0000000;
	124: instructionOdd = 32'h42001;
	125: instructionOdd = 32'hcbffff1;
	126: instructionOdd = 32'hf0080000;
	127: instructionOdd = 32'h400000;
	128: instructionOdd = 32'h4cbffffb;
	129: instructionOdd = 32'hf0080000;
	130: instructionOdd = 32'h87c40000;
	131: instructionOdd = 32'h2842080;
	132: instructionOdd = 32'h2022036;
	133: instructionOdd = 32'h40078;
	134: instructionOdd = 32'hf0080000;
	135: instructionOdd = 32'h87c40000;
	136: instructionOdd = 32'h2842080;
	137: instructionOdd = 32'h2022036;
	138: instructionOdd = 32'h87c40000;
	139: instructionOdd = 32'h2c22081;
	140: instructionOdd = 32'h2c60085;
	141: instructionOdd = 32'hf0000000;
	142: instructionOdd = 32'h20001;
	143: instructionOdd = 32'hc80000c;
	144: instructionOdd = 32'h2842189;
	145: instructionOdd = 32'h2022260;
	146: instructionOdd = 32'h87c40000;
	147: instructionOdd = 32'h2842082;
	148: instructionOdd = 32'h2021134;
	149: instructionOdd = 32'h87c40000;
	150: instructionOdd = 32'h20001;
	151: instructionOdd = 32'h2c22085;
	152: instructionOdd = 32'h2c22085;
	153: instructionOdd = 32'h2aff105;
	154: instructionOdd = 32'h2b3f107;
	155: instructionOdd = 32'h293f102;
	156: instructionOdd = 32'h2409028;
	157: instructionOdd = 32'h400000;
	158: instructionOdd = 32'h293f100;
	159: instructionOdd = 32'h20000;
	160: instructionOdd = 32'h3ff024;
	161: instructionOdd = 32'h7ff040;
	162: instructionOdd = 32'h2c5f487;
	163: instructionOdd = 32'h20000;
	164: instructionOdd = 32'h2c5fe0f;
	165: instructionOdd = 32'h2c5f486;
	166: instructionOdd = 32'h2c5f485;
	167: instructionOdd = 32'h2c5fb09;
	168: instructionOdd = 32'h2c5fc0b;
	169: instructionOdd = 32'h2c5fd0d;
	170: instructionOdd = 32'h20000;
	171: instructionOdd = 32'h20004;
	172: instructionOdd = 32'h2d41100;
	173: instructionOdd = 32'h20000;
	174: instructionOdd = 32'h400000;
	175: instructionOdd = 32'h2c42080;
	176: instructionOdd = 32'h2021134;
	177: instructionOdd = 32'h87c40000;
	178: instructionOdd = 32'h2c42080;
	179: instructionOdd = 32'h80000;
	180: instructionOdd = 32'h2c5f003;
	181: instructionOdd = 32'h340000;
	182: instructionOdd = 32'h2c5f002;
	183: instructionOdd = 32'h2c5f001;
	184: instructionOdd = 32'h20408;
	185: instructionOdd = 32'h420001;
	186: instructionOdd = 32'h40000;
	187: instructionOdd = 32'h381000;
	188: instructionOdd = 32'h2e3000;
	189: instructionOdd = 32'h87c20000;
	190: instructionOdd = 32'h2c21d80;
	191: instructionOdd = 32'h440001;
	192: instructionOdd = 32'hcfffff6;
	193: instructionOdd = 32'h60000;
	194: instructionOdd = 32'h2022b34;
	195: instructionOdd = 32'hc57008;
	196: instructionOdd = 32'h2061106;
	197: instructionOdd = 32'h5c004;
	198: instructionOdd = 32'hc800025;
	199: instructionOdd = 32'h60008;
	200: instructionOdd = 32'h2024036;
	201: instructionOdd = 32'hedb88320;
	202: instructionOdd = 32'h9044001;
	203: instructionOdd = 32'h463001;
	204: instructionOdd = 32'hcbffff7;
	205: instructionOdd = 32'h206300b;
	206: instructionOdd = 32'h28bf103;
	207: instructionOdd = 32'h20a1286;
	208: instructionOdd = 32'h2021db4;
	209: instructionOdd = 32'h289f102;
	210: instructionOdd = 32'h2023261;
	211: instructionOdd = 32'h20004;
	212: instructionOdd = 32'hc800018;
	213: instructionOdd = 32'hf0008010;
	214: instructionOdd = 32'h25000;
	215: instructionOdd = 32'h4c00012;
	216: instructionOdd = 32'h2c5f284;
	217: instructionOdd = 32'h59000;
	218: instructionOdd = 32'h2035c00;
	219: instructionOdd = 32'hfffffffc;
	220: instructionOdd = 32'h4c0000c;
	221: instructionOdd = 32'h400000;
	222: instructionOdd = 32'h4800004;
	223: instructionOdd = 32'h4800002;
	224: instructionOdd = 32'h283f101;
	225: instructionOdd = 32'h37b001;
	226: instructionOdd = 32'h2023230;
	227: instructionOdd = 32'h20220c7;
	228: instructionOdd = 32'h64003;
	229: instructionOdd = 32'hfffffffc;
	230: instructionOdd = 32'hcc0000a;
	231: instructionOdd = 32'h2c5f202;
	232: instructionOdd = 32'h63004;
	233: instructionOdd = 32'hcfffffd;
	234: instructionOdd = 32'hfffffffc;
	235: instructionOdd = 32'h360002;
	236: instructionOdd = 32'h287f100;
	237: instructionOdd = 32'h63001;
	238: instructionOdd = 32'h2c5f202;
	239: instructionOdd = 32'h1c75003;
	240: instructionOdd = 32'h80a0000;
	241: instructionOdd = 32'h2c5f081;
	242: instructionOdd = 32'h3c003;
	243: instructionOdd = 32'hcffff90;
	244: instructionOdd = 32'h3c000;
	245: instructionOdd = 32'hf0080000;
	246: instructionOdd = 32'h400000;
	247: instructionOdd = 32'h4cbffffb;
	248: instructionOdd = 32'h1c410ff;
	249: instructionOdd = 32'hf0080000;
	250: instructionOdd = 32'hcc0000c;
	251: instructionOdd = 32'h20000;
	252: instructionOdd = 32'h285f104;
	253: instructionOdd = 32'h2021131;
	254: instructionOdd = 32'h20000;
	255: instructionOdd = 32'h283f101;
	256: instructionOdd = 32'h2adf109;
	257: instructionOdd = 32'h2b1f10b;
	258: instructionOdd = 32'h2b5f10d;
	259: instructionOdd = 32'h2b9f10f;
	260: instructionOdd = 32'h2abf108;
	261: instructionOdd = 32'h293f106;
	262: instructionOdd = 32'h2409027;
	263: instructionOdd = 32'h6400000;
	264: instructionOdd = 32'h2409020;
	265: instructionOdd = 32'h1a4;
	266: instructionOdd = 32'h20000;
	267: instructionOdd = 32'h20404;
	268: instructionOdd = 32'h2842100;
	269: instructionOdd = 32'h20220b1;
	270: instructionOdd = 32'h87c40000;
	271: instructionOdd = 32'h2822100;
	272: instructionOdd = 32'h1021001;
	273: instructionOdd = 32'hcc00012;
	274: instructionOdd = 32'h2c42080;
	275: instructionOdd = 32'hf0080000;
	276: instructionOdd = 32'h400000;
	277: instructionOdd = 32'h2021060;
	278: instructionOdd = 32'h87c20000;
	279: instructionOdd = 32'h2821081;
	280: instructionOdd = 32'h20408;
	281: instructionOdd = 32'hff00;
	282: instructionOdd = 32'h1c41001;
	283: instructionOdd = 32'hf0080000;
	284: instructionOdd = 32'h400000;
	285: instructionOdd = 32'h2021060;
	286: instructionOdd = 32'h2022060;
	287: instructionOdd = 32'hf0080000;
	288: instructionOdd = 32'h2821081;
	289: instructionOdd = 32'h87c40000;
	290: instructionOdd = 32'h2862100;
	291: instructionOdd = 32'h87c83000;
	292: instructionOdd = 32'h2d44080;
	293: instructionOdd = 32'h4c00026;
	294: instructionOdd = 32'h2c42080;
	295: instructionOdd = 32'hf0080000;
	296: instructionOdd = 32'h400000;
	297: instructionOdd = 32'h2022060;
	298: instructionOdd = 32'h87c40000;
	299: instructionOdd = 32'h2862081;
	300: instructionOdd = 32'hc43002;
	301: instructionOdd = 32'h2022086;
	302: instructionOdd = 32'h20000;
	303: instructionOdd = 32'h1c6303f;
	304: instructionOdd = 32'h63002;
	305: instructionOdd = 32'h87c84000;
	306: instructionOdd = 32'h2884900;
	307: instructionOdd = 32'h20004;
	308: instructionOdd = 32'h20211b2;
	309: instructionOdd = 32'hcfffff7;
	310: instructionOdd = 32'h1c423ff;
	311: instructionOdd = 32'h20000;
	312: instructionOdd = 32'h87c40000;
	313: instructionOdd = 32'h2862100;
	314: instructionOdd = 32'h87c23000;
	315: instructionOdd = 32'h63001;
	316: instructionOdd = 32'h6400000;
	317: instructionOdd = 32'h2c42180;
	318: instructionOdd = 32'h0;
	319: instructionOdd = 32'h0;
	320: instructionOdd = 32'h0;
	321: instructionOdd = 32'h0;
	322: instructionOdd = 32'h0;
	323: instructionOdd = 32'h0;
	324: instructionOdd = 32'h0;
	325: instructionOdd = 32'h0;
	326: instructionOdd = 32'h0;
	327: instructionOdd = 32'h0;
	328: instructionOdd = 32'h0;
	329: instructionOdd = 32'h0;
	330: instructionOdd = 32'h0;
	331: instructionOdd = 32'h0;
	332: instructionOdd = 32'h0;
	333: instructionOdd = 32'h0;
	334: instructionOdd = 32'h0;
	335: instructionOdd = 32'h0;
	336: instructionOdd = 32'h0;
	337: instructionOdd = 32'h0;
	338: instructionOdd = 32'h0;
	339: instructionOdd = 32'h0;
	340: instructionOdd = 32'h0;
	341: instructionOdd = 32'h0;
	342: instructionOdd = 32'h0;
	343: instructionOdd = 32'h0;
	344: instructionOdd = 32'h0;
	345: instructionOdd = 32'h0;
	346: instructionOdd = 32'h0;
	347: instructionOdd = 32'h0;
	348: instructionOdd = 32'h0;
	349: instructionOdd = 32'h0;
	350: instructionOdd = 32'h0;
	351: instructionOdd = 32'h0;
	352: instructionOdd = 32'h0;
	353: instructionOdd = 32'h0;
	354: instructionOdd = 32'h0;
	355: instructionOdd = 32'h0;
	356: instructionOdd = 32'h0;
	357: instructionOdd = 32'h0;
	358: instructionOdd = 32'h0;
	359: instructionOdd = 32'h0;
	360: instructionOdd = 32'h0;
	361: instructionOdd = 32'h0;
	362: instructionOdd = 32'h0;
	363: instructionOdd = 32'h0;
	364: instructionOdd = 32'h0;
	365: instructionOdd = 32'h0;
	366: instructionOdd = 32'h0;
	367: instructionOdd = 32'h0;
	368: instructionOdd = 32'h0;
	369: instructionOdd = 32'h0;
	370: instructionOdd = 32'h0;
	371: instructionOdd = 32'h0;
	372: instructionOdd = 32'h0;
	373: instructionOdd = 32'h0;
	374: instructionOdd = 32'h0;
	375: instructionOdd = 32'h0;
	376: instructionOdd = 32'h0;
	377: instructionOdd = 32'h0;
	378: instructionOdd = 32'h0;
	379: instructionOdd = 32'h0;
	380: instructionOdd = 32'h0;
	381: instructionOdd = 32'h0;
	382: instructionOdd = 32'h0;
	383: instructionOdd = 32'h0;
	384: instructionOdd = 32'h0;
	385: instructionOdd = 32'h0;
	386: instructionOdd = 32'h0;
	387: instructionOdd = 32'h0;
	388: instructionOdd = 32'h0;
	389: instructionOdd = 32'h0;
	390: instructionOdd = 32'h0;
	391: instructionOdd = 32'h0;
	392: instructionOdd = 32'h0;
	393: instructionOdd = 32'h0;
	394: instructionOdd = 32'h0;
	395: instructionOdd = 32'h0;
	396: instructionOdd = 32'h0;
	397: instructionOdd = 32'h0;
	398: instructionOdd = 32'h0;
	399: instructionOdd = 32'h0;
	400: instructionOdd = 32'h0;
	401: instructionOdd = 32'h0;
	402: instructionOdd = 32'h0;
	403: instructionOdd = 32'h0;
	404: instructionOdd = 32'h0;
	405: instructionOdd = 32'h0;
	406: instructionOdd = 32'h0;
	407: instructionOdd = 32'h0;
	408: instructionOdd = 32'h0;
	409: instructionOdd = 32'h0;
	410: instructionOdd = 32'h0;
	411: instructionOdd = 32'h0;
	412: instructionOdd = 32'h0;
	413: instructionOdd = 32'h0;
	414: instructionOdd = 32'h0;
	415: instructionOdd = 32'h0;
	416: instructionOdd = 32'h0;
	417: instructionOdd = 32'h0;
	418: instructionOdd = 32'h0;
	419: instructionOdd = 32'h0;
	420: instructionOdd = 32'h0;
	421: instructionOdd = 32'h0;
	422: instructionOdd = 32'h0;
	423: instructionOdd = 32'h0;
	424: instructionOdd = 32'h0;
	425: instructionOdd = 32'h0;
	426: instructionOdd = 32'h0;
	427: instructionOdd = 32'h0;
	428: instructionOdd = 32'h0;
	429: instructionOdd = 32'h0;
	430: instructionOdd = 32'h0;
	431: instructionOdd = 32'h0;
	432: instructionOdd = 32'h0;
	433: instructionOdd = 32'h0;
	434: instructionOdd = 32'h0;
	435: instructionOdd = 32'h0;
	436: instructionOdd = 32'h0;
	437: instructionOdd = 32'h0;
	438: instructionOdd = 32'h0;
	439: instructionOdd = 32'h0;
	440: instructionOdd = 32'h0;
	441: instructionOdd = 32'h0;
	442: instructionOdd = 32'h0;
	443: instructionOdd = 32'h0;
	444: instructionOdd = 32'h0;
	445: instructionOdd = 32'h0;
	446: instructionOdd = 32'h0;
	447: instructionOdd = 32'h0;
	448: instructionOdd = 32'h0;
	449: instructionOdd = 32'h0;
	450: instructionOdd = 32'h0;
	451: instructionOdd = 32'h0;
	452: instructionOdd = 32'h0;
	453: instructionOdd = 32'h0;
	454: instructionOdd = 32'h0;
	455: instructionOdd = 32'h0;
	456: instructionOdd = 32'h0;
	457: instructionOdd = 32'h0;
	458: instructionOdd = 32'h0;
	459: instructionOdd = 32'h0;
	460: instructionOdd = 32'h0;
	461: instructionOdd = 32'h0;
	462: instructionOdd = 32'h0;
	463: instructionOdd = 32'h0;
	464: instructionOdd = 32'h0;
	465: instructionOdd = 32'h0;
	466: instructionOdd = 32'h0;
	467: instructionOdd = 32'h0;
	468: instructionOdd = 32'h0;
	469: instructionOdd = 32'h0;
	470: instructionOdd = 32'h0;
	471: instructionOdd = 32'h0;
	472: instructionOdd = 32'h0;
	473: instructionOdd = 32'h0;
	474: instructionOdd = 32'h0;
	475: instructionOdd = 32'h0;
	476: instructionOdd = 32'h0;
	477: instructionOdd = 32'h0;
	478: instructionOdd = 32'h0;
	479: instructionOdd = 32'h0;
	480: instructionOdd = 32'h0;
	481: instructionOdd = 32'h0;
	482: instructionOdd = 32'h0;
	483: instructionOdd = 32'h0;
	484: instructionOdd = 32'h0;
	485: instructionOdd = 32'h0;
	486: instructionOdd = 32'h0;
	487: instructionOdd = 32'h0;
	488: instructionOdd = 32'h0;
	489: instructionOdd = 32'h0;
	490: instructionOdd = 32'h0;
	491: instructionOdd = 32'h0;
	492: instructionOdd = 32'h0;
	493: instructionOdd = 32'h0;
	494: instructionOdd = 32'h0;
	495: instructionOdd = 32'h0;
	496: instructionOdd = 32'h0;
	497: instructionOdd = 32'h0;
	498: instructionOdd = 32'h0;
	499: instructionOdd = 32'h0;
	500: instructionOdd = 32'h0;
	501: instructionOdd = 32'h0;
	502: instructionOdd = 32'h0;
	503: instructionOdd = 32'h0;
	504: instructionOdd = 32'h0;
	505: instructionOdd = 32'h0;
	506: instructionOdd = 32'h0;
	507: instructionOdd = 32'h0;
	508: instructionOdd = 32'h0;
	509: instructionOdd = 32'h0;
	510: instructionOdd = 32'h0;
	511: instructionOdd = 32'h0;
	512: instructionOdd = 32'h0;
	513: instructionOdd = 32'h0;
	514: instructionOdd = 32'h0;
	515: instructionOdd = 32'h0;
	516: instructionOdd = 32'h0;
	517: instructionOdd = 32'h0;
	518: instructionOdd = 32'h0;
	519: instructionOdd = 32'h0;
	520: instructionOdd = 32'h0;
	521: instructionOdd = 32'h0;
	522: instructionOdd = 32'h0;
	523: instructionOdd = 32'h0;
	524: instructionOdd = 32'h0;
	525: instructionOdd = 32'h0;
	526: instructionOdd = 32'h0;
	527: instructionOdd = 32'h0;
	528: instructionOdd = 32'h0;
	529: instructionOdd = 32'h0;
	530: instructionOdd = 32'h0;
	531: instructionOdd = 32'h0;
	532: instructionOdd = 32'h0;
	533: instructionOdd = 32'h0;
	534: instructionOdd = 32'h0;
	535: instructionOdd = 32'h0;
	536: instructionOdd = 32'h0;
	537: instructionOdd = 32'h0;
	538: instructionOdd = 32'h0;
	539: instructionOdd = 32'h0;
	540: instructionOdd = 32'h0;
	541: instructionOdd = 32'h0;
	542: instructionOdd = 32'h0;
	543: instructionOdd = 32'h0;
	544: instructionOdd = 32'h0;
	545: instructionOdd = 32'h0;
	546: instructionOdd = 32'h0;
	547: instructionOdd = 32'h0;
	548: instructionOdd = 32'h0;
	549: instructionOdd = 32'h0;
	550: instructionOdd = 32'h0;
	551: instructionOdd = 32'h0;
	552: instructionOdd = 32'h0;
	553: instructionOdd = 32'h0;
	554: instructionOdd = 32'h0;
	555: instructionOdd = 32'h0;
	556: instructionOdd = 32'h0;
	557: instructionOdd = 32'h0;
	558: instructionOdd = 32'h0;
	559: instructionOdd = 32'h0;
	560: instructionOdd = 32'h0;
	561: instructionOdd = 32'h0;
	562: instructionOdd = 32'h0;
	563: instructionOdd = 32'h0;
	564: instructionOdd = 32'h0;
	565: instructionOdd = 32'h0;
	566: instructionOdd = 32'h0;
	567: instructionOdd = 32'h0;
	568: instructionOdd = 32'h0;
	569: instructionOdd = 32'h0;
	570: instructionOdd = 32'h0;
	571: instructionOdd = 32'h0;
	572: instructionOdd = 32'h0;
	573: instructionOdd = 32'h0;
	574: instructionOdd = 32'h0;
	575: instructionOdd = 32'h0;
	576: instructionOdd = 32'h0;
	577: instructionOdd = 32'h0;
	578: instructionOdd = 32'h0;
	579: instructionOdd = 32'h0;
	580: instructionOdd = 32'h0;
	581: instructionOdd = 32'h0;
	582: instructionOdd = 32'h0;
	583: instructionOdd = 32'h0;
	584: instructionOdd = 32'h0;
	585: instructionOdd = 32'h0;
	586: instructionOdd = 32'h0;
	587: instructionOdd = 32'h0;
	588: instructionOdd = 32'h0;
	589: instructionOdd = 32'h0;
	590: instructionOdd = 32'h0;
	591: instructionOdd = 32'h0;
	592: instructionOdd = 32'h0;
	593: instructionOdd = 32'h0;
	594: instructionOdd = 32'h0;
	595: instructionOdd = 32'h0;
	596: instructionOdd = 32'h0;
	597: instructionOdd = 32'h0;
	598: instructionOdd = 32'h0;
	599: instructionOdd = 32'h0;
	600: instructionOdd = 32'h0;
	601: instructionOdd = 32'h0;
	602: instructionOdd = 32'h0;
	603: instructionOdd = 32'h0;
	604: instructionOdd = 32'h0;
	605: instructionOdd = 32'h0;
	606: instructionOdd = 32'h0;
	607: instructionOdd = 32'h0;
	608: instructionOdd = 32'h0;
	609: instructionOdd = 32'h0;
	610: instructionOdd = 32'h0;
	611: instructionOdd = 32'h0;
	612: instructionOdd = 32'h0;
	613: instructionOdd = 32'h0;
	614: instructionOdd = 32'h0;
	615: instructionOdd = 32'h0;
	616: instructionOdd = 32'h0;
	617: instructionOdd = 32'h0;
	618: instructionOdd = 32'h0;
	619: instructionOdd = 32'h0;
	620: instructionOdd = 32'h0;
	621: instructionOdd = 32'h0;
	622: instructionOdd = 32'h0;
	623: instructionOdd = 32'h0;
	624: instructionOdd = 32'h0;
	625: instructionOdd = 32'h0;
	626: instructionOdd = 32'h0;
	627: instructionOdd = 32'h0;
	628: instructionOdd = 32'h0;
	629: instructionOdd = 32'h0;
	630: instructionOdd = 32'h0;
	631: instructionOdd = 32'h0;
	632: instructionOdd = 32'h0;
	633: instructionOdd = 32'h0;
	634: instructionOdd = 32'h0;
	635: instructionOdd = 32'h0;
	636: instructionOdd = 32'h0;
	637: instructionOdd = 32'h0;
	638: instructionOdd = 32'h0;
	639: instructionOdd = 32'h0;
	640: instructionOdd = 32'h0;
	641: instructionOdd = 32'h0;
	642: instructionOdd = 32'h0;
	643: instructionOdd = 32'h0;
	644: instructionOdd = 32'h0;
	645: instructionOdd = 32'h0;
	646: instructionOdd = 32'h0;
	647: instructionOdd = 32'h0;
	648: instructionOdd = 32'h0;
	649: instructionOdd = 32'h0;
	650: instructionOdd = 32'h0;
	651: instructionOdd = 32'h0;
	652: instructionOdd = 32'h0;
	653: instructionOdd = 32'h0;
	654: instructionOdd = 32'h0;
	655: instructionOdd = 32'h0;
	656: instructionOdd = 32'h0;
	657: instructionOdd = 32'h0;
	658: instructionOdd = 32'h0;
	659: instructionOdd = 32'h0;
	660: instructionOdd = 32'h0;
	661: instructionOdd = 32'h0;
	662: instructionOdd = 32'h0;
	663: instructionOdd = 32'h0;
	664: instructionOdd = 32'h0;
	665: instructionOdd = 32'h0;
	666: instructionOdd = 32'h0;
	667: instructionOdd = 32'h0;
	668: instructionOdd = 32'h0;
	669: instructionOdd = 32'h0;
	670: instructionOdd = 32'h0;
	671: instructionOdd = 32'h0;
	672: instructionOdd = 32'h0;
	673: instructionOdd = 32'h0;
	674: instructionOdd = 32'h0;
	675: instructionOdd = 32'h0;
	676: instructionOdd = 32'h0;
	677: instructionOdd = 32'h0;
	678: instructionOdd = 32'h0;
	679: instructionOdd = 32'h0;
	680: instructionOdd = 32'h0;
	681: instructionOdd = 32'h0;
	682: instructionOdd = 32'h0;
	683: instructionOdd = 32'h0;
	684: instructionOdd = 32'h0;
	685: instructionOdd = 32'h0;
	686: instructionOdd = 32'h0;
	687: instructionOdd = 32'h0;
	688: instructionOdd = 32'h0;
	689: instructionOdd = 32'h0;
	690: instructionOdd = 32'h0;
	691: instructionOdd = 32'h0;
	692: instructionOdd = 32'h0;
	693: instructionOdd = 32'h0;
	694: instructionOdd = 32'h0;
	695: instructionOdd = 32'h0;
	696: instructionOdd = 32'h0;
	697: instructionOdd = 32'h0;
	698: instructionOdd = 32'h0;
	699: instructionOdd = 32'h0;
	700: instructionOdd = 32'h0;
	701: instructionOdd = 32'h0;
	702: instructionOdd = 32'h0;
	703: instructionOdd = 32'h0;
	704: instructionOdd = 32'h0;
	705: instructionOdd = 32'h0;
	706: instructionOdd = 32'h0;
	707: instructionOdd = 32'h0;
	708: instructionOdd = 32'h0;
	709: instructionOdd = 32'h0;
	710: instructionOdd = 32'h0;
	711: instructionOdd = 32'h0;
	712: instructionOdd = 32'h0;
	713: instructionOdd = 32'h0;
	714: instructionOdd = 32'h0;
	715: instructionOdd = 32'h0;
	716: instructionOdd = 32'h0;
	717: instructionOdd = 32'h0;
	718: instructionOdd = 32'h0;
	719: instructionOdd = 32'h0;
	720: instructionOdd = 32'h0;
	721: instructionOdd = 32'h0;
	722: instructionOdd = 32'h0;
	723: instructionOdd = 32'h0;
	724: instructionOdd = 32'h0;
	725: instructionOdd = 32'h0;
	726: instructionOdd = 32'h0;
	727: instructionOdd = 32'h0;
	728: instructionOdd = 32'h0;
	729: instructionOdd = 32'h0;
	730: instructionOdd = 32'h0;
	731: instructionOdd = 32'h0;
	732: instructionOdd = 32'h0;
	733: instructionOdd = 32'h0;
	734: instructionOdd = 32'h0;
	735: instructionOdd = 32'h0;
	736: instructionOdd = 32'h0;
	737: instructionOdd = 32'h0;
	738: instructionOdd = 32'h0;
	739: instructionOdd = 32'h0;
	740: instructionOdd = 32'h0;
	741: instructionOdd = 32'h0;
	742: instructionOdd = 32'h0;
	743: instructionOdd = 32'h0;
	744: instructionOdd = 32'h0;
	745: instructionOdd = 32'h0;
	746: instructionOdd = 32'h0;
	747: instructionOdd = 32'h0;
	748: instructionOdd = 32'h0;
	749: instructionOdd = 32'h0;
	750: instructionOdd = 32'h0;
	751: instructionOdd = 32'h0;
	752: instructionOdd = 32'h0;
	753: instructionOdd = 32'h0;
	754: instructionOdd = 32'h0;
	755: instructionOdd = 32'h0;
	756: instructionOdd = 32'h0;
	757: instructionOdd = 32'h0;
	758: instructionOdd = 32'h0;
	759: instructionOdd = 32'h0;
	760: instructionOdd = 32'h0;
	761: instructionOdd = 32'h0;
	762: instructionOdd = 32'h0;
	763: instructionOdd = 32'h0;
	764: instructionOdd = 32'h0;
	765: instructionOdd = 32'h0;
	766: instructionOdd = 32'h0;
	767: instructionOdd = 32'h0;
	768: instructionOdd = 32'h0;
	769: instructionOdd = 32'h0;
	770: instructionOdd = 32'h0;
	771: instructionOdd = 32'h0;
	772: instructionOdd = 32'h0;
	773: instructionOdd = 32'h0;
	774: instructionOdd = 32'h0;
	775: instructionOdd = 32'h0;
	776: instructionOdd = 32'h0;
	777: instructionOdd = 32'h0;
	778: instructionOdd = 32'h0;
	779: instructionOdd = 32'h0;
	780: instructionOdd = 32'h0;
	781: instructionOdd = 32'h0;
	782: instructionOdd = 32'h0;
	783: instructionOdd = 32'h0;
	784: instructionOdd = 32'h0;
	785: instructionOdd = 32'h0;
	786: instructionOdd = 32'h0;
	787: instructionOdd = 32'h0;
	788: instructionOdd = 32'h0;
	789: instructionOdd = 32'h0;
	790: instructionOdd = 32'h0;
	791: instructionOdd = 32'h0;
	792: instructionOdd = 32'h0;
	793: instructionOdd = 32'h0;
	794: instructionOdd = 32'h0;
	795: instructionOdd = 32'h0;
	796: instructionOdd = 32'h0;
	797: instructionOdd = 32'h0;
	798: instructionOdd = 32'h0;
	799: instructionOdd = 32'h0;
	800: instructionOdd = 32'h0;
	801: instructionOdd = 32'h0;
	802: instructionOdd = 32'h0;
	803: instructionOdd = 32'h0;
	804: instructionOdd = 32'h0;
	805: instructionOdd = 32'h0;
	806: instructionOdd = 32'h0;
	807: instructionOdd = 32'h0;
	808: instructionOdd = 32'h0;
	809: instructionOdd = 32'h0;
	810: instructionOdd = 32'h0;
	811: instructionOdd = 32'h0;
	812: instructionOdd = 32'h0;
	813: instructionOdd = 32'h0;
	814: instructionOdd = 32'h0;
	815: instructionOdd = 32'h0;
	816: instructionOdd = 32'h0;
	817: instructionOdd = 32'h0;
	818: instructionOdd = 32'h0;
	819: instructionOdd = 32'h0;
	820: instructionOdd = 32'h0;
	821: instructionOdd = 32'h0;
	822: instructionOdd = 32'h0;
	823: instructionOdd = 32'h0;
	824: instructionOdd = 32'h0;
	825: instructionOdd = 32'h0;
	826: instructionOdd = 32'h0;
	827: instructionOdd = 32'h0;
	828: instructionOdd = 32'h0;
	829: instructionOdd = 32'h0;
	830: instructionOdd = 32'h0;
	831: instructionOdd = 32'h0;
	832: instructionOdd = 32'h0;
	833: instructionOdd = 32'h0;
	834: instructionOdd = 32'h0;
	835: instructionOdd = 32'h0;
	836: instructionOdd = 32'h0;
	837: instructionOdd = 32'h0;
	838: instructionOdd = 32'h0;
	839: instructionOdd = 32'h0;
	840: instructionOdd = 32'h0;
	841: instructionOdd = 32'h0;
	842: instructionOdd = 32'h0;
	843: instructionOdd = 32'h0;
	844: instructionOdd = 32'h0;
	845: instructionOdd = 32'h0;
	846: instructionOdd = 32'h0;
	847: instructionOdd = 32'h0;
	848: instructionOdd = 32'h0;
	849: instructionOdd = 32'h0;
	850: instructionOdd = 32'h0;
	851: instructionOdd = 32'h0;
	852: instructionOdd = 32'h0;
	853: instructionOdd = 32'h0;
	854: instructionOdd = 32'h0;
	855: instructionOdd = 32'h0;
	856: instructionOdd = 32'h0;
	857: instructionOdd = 32'h0;
	858: instructionOdd = 32'h0;
	859: instructionOdd = 32'h0;
	860: instructionOdd = 32'h0;
	861: instructionOdd = 32'h0;
	862: instructionOdd = 32'h0;
	863: instructionOdd = 32'h0;
	864: instructionOdd = 32'h0;
	865: instructionOdd = 32'h0;
	866: instructionOdd = 32'h0;
	867: instructionOdd = 32'h0;
	868: instructionOdd = 32'h0;
	869: instructionOdd = 32'h0;
	870: instructionOdd = 32'h0;
	871: instructionOdd = 32'h0;
	872: instructionOdd = 32'h0;
	873: instructionOdd = 32'h0;
	874: instructionOdd = 32'h0;
	875: instructionOdd = 32'h0;
	876: instructionOdd = 32'h0;
	877: instructionOdd = 32'h0;
	878: instructionOdd = 32'h0;
	879: instructionOdd = 32'h0;
	880: instructionOdd = 32'h0;
	881: instructionOdd = 32'h0;
	882: instructionOdd = 32'h0;
	883: instructionOdd = 32'h0;
	884: instructionOdd = 32'h0;
	885: instructionOdd = 32'h0;
	886: instructionOdd = 32'h0;
	887: instructionOdd = 32'h0;
	888: instructionOdd = 32'h0;
	889: instructionOdd = 32'h0;
	890: instructionOdd = 32'h0;
	891: instructionOdd = 32'h0;
	892: instructionOdd = 32'h0;
	893: instructionOdd = 32'h0;
	894: instructionOdd = 32'h0;
	895: instructionOdd = 32'h0;
	896: instructionOdd = 32'h0;
	897: instructionOdd = 32'h0;
	898: instructionOdd = 32'h0;
	899: instructionOdd = 32'h0;
	900: instructionOdd = 32'h0;
	901: instructionOdd = 32'h0;
	902: instructionOdd = 32'h0;
	903: instructionOdd = 32'h0;
	904: instructionOdd = 32'h0;
	905: instructionOdd = 32'h0;
	906: instructionOdd = 32'h0;
	907: instructionOdd = 32'h0;
	908: instructionOdd = 32'h0;
	909: instructionOdd = 32'h0;
	910: instructionOdd = 32'h0;
	911: instructionOdd = 32'h0;
	912: instructionOdd = 32'h0;
	913: instructionOdd = 32'h0;
	914: instructionOdd = 32'h0;
	915: instructionOdd = 32'h0;
	916: instructionOdd = 32'h0;
	917: instructionOdd = 32'h0;
	918: instructionOdd = 32'h0;
	919: instructionOdd = 32'h0;
	920: instructionOdd = 32'h0;
	921: instructionOdd = 32'h0;
	922: instructionOdd = 32'h0;
	923: instructionOdd = 32'h0;
	924: instructionOdd = 32'h0;
	925: instructionOdd = 32'h0;
	926: instructionOdd = 32'h0;
	927: instructionOdd = 32'h0;
	928: instructionOdd = 32'h0;
	929: instructionOdd = 32'h0;
	930: instructionOdd = 32'h0;
	931: instructionOdd = 32'h0;
	932: instructionOdd = 32'h0;
	933: instructionOdd = 32'h0;
	934: instructionOdd = 32'h0;
	935: instructionOdd = 32'h0;
	936: instructionOdd = 32'h0;
	937: instructionOdd = 32'h0;
	938: instructionOdd = 32'h0;
	939: instructionOdd = 32'h0;
	940: instructionOdd = 32'h0;
	941: instructionOdd = 32'h0;
	942: instructionOdd = 32'h0;
	943: instructionOdd = 32'h0;
	944: instructionOdd = 32'h0;
	945: instructionOdd = 32'h0;
	946: instructionOdd = 32'h0;
	947: instructionOdd = 32'h0;
	948: instructionOdd = 32'h0;
	949: instructionOdd = 32'h0;
	950: instructionOdd = 32'h0;
	951: instructionOdd = 32'h0;
	952: instructionOdd = 32'h0;
	953: instructionOdd = 32'h0;
	954: instructionOdd = 32'h0;
	955: instructionOdd = 32'h0;
	956: instructionOdd = 32'h0;
	957: instructionOdd = 32'h0;
	958: instructionOdd = 32'h0;
	959: instructionOdd = 32'h0;
	960: instructionOdd = 32'h0;
	961: instructionOdd = 32'h0;
	962: instructionOdd = 32'h0;
	963: instructionOdd = 32'h0;
	964: instructionOdd = 32'h0;
	965: instructionOdd = 32'h0;
	966: instructionOdd = 32'h0;
	967: instructionOdd = 32'h0;
	968: instructionOdd = 32'h0;
	969: instructionOdd = 32'h0;
	970: instructionOdd = 32'h0;
	971: instructionOdd = 32'h0;
	972: instructionOdd = 32'h0;
	973: instructionOdd = 32'h0;
	974: instructionOdd = 32'h0;
	975: instructionOdd = 32'h0;
	976: instructionOdd = 32'h0;
	977: instructionOdd = 32'h0;
	978: instructionOdd = 32'h0;
	979: instructionOdd = 32'h0;
	980: instructionOdd = 32'h0;
	981: instructionOdd = 32'h0;
	982: instructionOdd = 32'h0;
	983: instructionOdd = 32'h0;
	984: instructionOdd = 32'h0;
	985: instructionOdd = 32'h0;
	986: instructionOdd = 32'h0;
	987: instructionOdd = 32'h0;
	988: instructionOdd = 32'h0;
	989: instructionOdd = 32'h0;
	990: instructionOdd = 32'h0;
	991: instructionOdd = 32'h0;
	992: instructionOdd = 32'h0;
	993: instructionOdd = 32'h0;
	994: instructionOdd = 32'h0;
	995: instructionOdd = 32'h0;
	996: instructionOdd = 32'h0;
	997: instructionOdd = 32'h0;
	998: instructionOdd = 32'h0;
	999: instructionOdd = 32'h0;
	1000: instructionOdd = 32'h0;
	1001: instructionOdd = 32'h0;
	1002: instructionOdd = 32'h0;
	1003: instructionOdd = 32'h0;
	1004: instructionOdd = 32'h0;
	1005: instructionOdd = 32'h0;
	1006: instructionOdd = 32'h0;
	1007: instructionOdd = 32'h0;
	1008: instructionOdd = 32'h0;
	1009: instructionOdd = 32'h0;
	1010: instructionOdd = 32'h0;
	1011: instructionOdd = 32'h0;
	1012: instructionOdd = 32'h0;
	1013: instructionOdd = 32'h0;
	1014: instructionOdd = 32'h0;
	1015: instructionOdd = 32'h0;
	1016: instructionOdd = 32'h0;
	1017: instructionOdd = 32'h0;
	1018: instructionOdd = 32'h0;
	1019: instructionOdd = 32'h0;
	1020: instructionOdd = 32'h0;
	1021: instructionOdd = 32'h0;
	1022: instructionOdd = 32'h0;
	1023: instructionOdd = 32'h0;
	1024: instructionOdd = 32'h0;
	1025: instructionOdd = 32'h0;
	1026: instructionOdd = 32'h0;
	1027: instructionOdd = 32'h0;
	1028: instructionOdd = 32'h0;
	1029: instructionOdd = 32'h0;
	1030: instructionOdd = 32'h0;
	1031: instructionOdd = 32'h0;
	1032: instructionOdd = 32'h0;
	1033: instructionOdd = 32'h0;
	1034: instructionOdd = 32'h0;
	1035: instructionOdd = 32'h0;
	1036: instructionOdd = 32'h0;
	1037: instructionOdd = 32'h0;
	1038: instructionOdd = 32'h0;
	1039: instructionOdd = 32'h0;
	1040: instructionOdd = 32'h0;
	1041: instructionOdd = 32'h0;
	1042: instructionOdd = 32'h0;
	1043: instructionOdd = 32'h0;
	1044: instructionOdd = 32'h0;
	1045: instructionOdd = 32'h0;
	1046: instructionOdd = 32'h0;
	1047: instructionOdd = 32'h0;
	1048: instructionOdd = 32'h0;
	1049: instructionOdd = 32'h0;
	1050: instructionOdd = 32'h0;
	1051: instructionOdd = 32'h0;
	1052: instructionOdd = 32'h0;
	1053: instructionOdd = 32'h0;
	1054: instructionOdd = 32'h0;
	1055: instructionOdd = 32'h0;
	1056: instructionOdd = 32'h0;
	1057: instructionOdd = 32'h0;
	1058: instructionOdd = 32'h0;
	1059: instructionOdd = 32'h0;
	1060: instructionOdd = 32'h0;
	1061: instructionOdd = 32'h0;
	1062: instructionOdd = 32'h0;
	1063: instructionOdd = 32'h0;
	1064: instructionOdd = 32'h0;
	1065: instructionOdd = 32'h0;
	1066: instructionOdd = 32'h0;
	1067: instructionOdd = 32'h0;
	1068: instructionOdd = 32'h0;
	1069: instructionOdd = 32'h0;
	1070: instructionOdd = 32'h0;
	1071: instructionOdd = 32'h0;
	1072: instructionOdd = 32'h0;
	1073: instructionOdd = 32'h0;
	1074: instructionOdd = 32'h0;
	1075: instructionOdd = 32'h0;
	1076: instructionOdd = 32'h0;
	1077: instructionOdd = 32'h0;
	1078: instructionOdd = 32'h0;
	1079: instructionOdd = 32'h0;
	1080: instructionOdd = 32'h0;
	1081: instructionOdd = 32'h0;
	1082: instructionOdd = 32'h0;
	1083: instructionOdd = 32'h0;
	1084: instructionOdd = 32'h0;
	1085: instructionOdd = 32'h0;
	1086: instructionOdd = 32'h0;
	1087: instructionOdd = 32'h0;
	1088: instructionOdd = 32'h0;
	1089: instructionOdd = 32'h0;
	1090: instructionOdd = 32'h0;
	1091: instructionOdd = 32'h0;
	1092: instructionOdd = 32'h0;
	1093: instructionOdd = 32'h0;
	1094: instructionOdd = 32'h0;
	1095: instructionOdd = 32'h0;
	1096: instructionOdd = 32'h0;
	1097: instructionOdd = 32'h0;
	1098: instructionOdd = 32'h0;
	1099: instructionOdd = 32'h0;
	1100: instructionOdd = 32'h0;
	1101: instructionOdd = 32'h0;
	1102: instructionOdd = 32'h0;
	1103: instructionOdd = 32'h0;
	1104: instructionOdd = 32'h0;
	1105: instructionOdd = 32'h0;
	1106: instructionOdd = 32'h0;
	1107: instructionOdd = 32'h0;
	1108: instructionOdd = 32'h0;
	1109: instructionOdd = 32'h0;
	1110: instructionOdd = 32'h0;
	1111: instructionOdd = 32'h0;
	1112: instructionOdd = 32'h0;
	1113: instructionOdd = 32'h0;
	1114: instructionOdd = 32'h0;
	1115: instructionOdd = 32'h0;
	1116: instructionOdd = 32'h0;
	1117: instructionOdd = 32'h0;
	1118: instructionOdd = 32'h0;
	1119: instructionOdd = 32'h0;
	1120: instructionOdd = 32'h0;
	1121: instructionOdd = 32'h0;
	1122: instructionOdd = 32'h0;
	1123: instructionOdd = 32'h0;
	1124: instructionOdd = 32'h0;
	1125: instructionOdd = 32'h0;
	1126: instructionOdd = 32'h0;
	1127: instructionOdd = 32'h0;
	1128: instructionOdd = 32'h0;
	1129: instructionOdd = 32'h0;
	1130: instructionOdd = 32'h0;
	1131: instructionOdd = 32'h0;
	1132: instructionOdd = 32'h0;
	1133: instructionOdd = 32'h0;
	1134: instructionOdd = 32'h0;
	1135: instructionOdd = 32'h0;
	1136: instructionOdd = 32'h0;
	1137: instructionOdd = 32'h0;
	1138: instructionOdd = 32'h0;
	1139: instructionOdd = 32'h0;
	1140: instructionOdd = 32'h0;
	1141: instructionOdd = 32'h0;
	1142: instructionOdd = 32'h0;
	1143: instructionOdd = 32'h0;
	1144: instructionOdd = 32'h0;
	1145: instructionOdd = 32'h0;
	1146: instructionOdd = 32'h0;
	1147: instructionOdd = 32'h0;
	1148: instructionOdd = 32'h0;
	1149: instructionOdd = 32'h0;
	1150: instructionOdd = 32'h0;
	1151: instructionOdd = 32'h0;
	1152: instructionOdd = 32'h0;
	1153: instructionOdd = 32'h0;
	1154: instructionOdd = 32'h0;
	1155: instructionOdd = 32'h0;
	1156: instructionOdd = 32'h0;
	1157: instructionOdd = 32'h0;
	1158: instructionOdd = 32'h0;
	1159: instructionOdd = 32'h0;
	1160: instructionOdd = 32'h0;
	1161: instructionOdd = 32'h0;
	1162: instructionOdd = 32'h0;
	1163: instructionOdd = 32'h0;
	1164: instructionOdd = 32'h0;
	1165: instructionOdd = 32'h0;
	1166: instructionOdd = 32'h0;
	1167: instructionOdd = 32'h0;
	1168: instructionOdd = 32'h0;
	1169: instructionOdd = 32'h0;
	1170: instructionOdd = 32'h0;
	1171: instructionOdd = 32'h0;
	1172: instructionOdd = 32'h0;
	1173: instructionOdd = 32'h0;
	1174: instructionOdd = 32'h0;
	1175: instructionOdd = 32'h0;
	1176: instructionOdd = 32'h0;
	1177: instructionOdd = 32'h0;
	1178: instructionOdd = 32'h0;
	1179: instructionOdd = 32'h0;
	1180: instructionOdd = 32'h0;
	1181: instructionOdd = 32'h0;
	1182: instructionOdd = 32'h0;
	1183: instructionOdd = 32'h0;
	1184: instructionOdd = 32'h0;
	1185: instructionOdd = 32'h0;
	1186: instructionOdd = 32'h0;
	1187: instructionOdd = 32'h0;
	1188: instructionOdd = 32'h0;
	1189: instructionOdd = 32'h0;
	1190: instructionOdd = 32'h0;
	1191: instructionOdd = 32'h0;
	1192: instructionOdd = 32'h0;
	1193: instructionOdd = 32'h0;
	1194: instructionOdd = 32'h0;
	1195: instructionOdd = 32'h0;
	1196: instructionOdd = 32'h0;
	1197: instructionOdd = 32'h0;
	1198: instructionOdd = 32'h0;
	1199: instructionOdd = 32'h0;
	1200: instructionOdd = 32'h0;
	1201: instructionOdd = 32'h0;
	1202: instructionOdd = 32'h0;
	1203: instructionOdd = 32'h0;
	1204: instructionOdd = 32'h0;
	1205: instructionOdd = 32'h0;
	1206: instructionOdd = 32'h0;
	1207: instructionOdd = 32'h0;
	1208: instructionOdd = 32'h0;
	1209: instructionOdd = 32'h0;
	1210: instructionOdd = 32'h0;
	1211: instructionOdd = 32'h0;
	1212: instructionOdd = 32'h0;
	1213: instructionOdd = 32'h0;
	1214: instructionOdd = 32'h0;
	1215: instructionOdd = 32'h0;
	1216: instructionOdd = 32'h0;
	1217: instructionOdd = 32'h0;
	1218: instructionOdd = 32'h0;
	1219: instructionOdd = 32'h0;
	1220: instructionOdd = 32'h0;
	1221: instructionOdd = 32'h0;
	1222: instructionOdd = 32'h0;
	1223: instructionOdd = 32'h0;
	1224: instructionOdd = 32'h0;
	1225: instructionOdd = 32'h0;
	1226: instructionOdd = 32'h0;
	1227: instructionOdd = 32'h0;
	1228: instructionOdd = 32'h0;
	1229: instructionOdd = 32'h0;
	1230: instructionOdd = 32'h0;
	1231: instructionOdd = 32'h0;
	1232: instructionOdd = 32'h0;
	1233: instructionOdd = 32'h0;
	1234: instructionOdd = 32'h0;
	1235: instructionOdd = 32'h0;
	1236: instructionOdd = 32'h0;
	1237: instructionOdd = 32'h0;
	1238: instructionOdd = 32'h0;
	1239: instructionOdd = 32'h0;
	1240: instructionOdd = 32'h0;
	1241: instructionOdd = 32'h0;
	1242: instructionOdd = 32'h0;
	1243: instructionOdd = 32'h0;
	1244: instructionOdd = 32'h0;
	1245: instructionOdd = 32'h0;
	1246: instructionOdd = 32'h0;
	1247: instructionOdd = 32'h0;
	1248: instructionOdd = 32'h0;
	1249: instructionOdd = 32'h0;
	1250: instructionOdd = 32'h0;
	1251: instructionOdd = 32'h0;
	1252: instructionOdd = 32'h0;
	1253: instructionOdd = 32'h0;
	1254: instructionOdd = 32'h0;
	1255: instructionOdd = 32'h0;
	1256: instructionOdd = 32'h0;
	1257: instructionOdd = 32'h0;
	1258: instructionOdd = 32'h0;
	1259: instructionOdd = 32'h0;
	1260: instructionOdd = 32'h0;
	1261: instructionOdd = 32'h0;
	1262: instructionOdd = 32'h0;
	1263: instructionOdd = 32'h0;
	1264: instructionOdd = 32'h0;
	1265: instructionOdd = 32'h0;
	1266: instructionOdd = 32'h0;
	1267: instructionOdd = 32'h0;
	1268: instructionOdd = 32'h0;
	1269: instructionOdd = 32'h0;
	1270: instructionOdd = 32'h0;
	1271: instructionOdd = 32'h0;
	1272: instructionOdd = 32'h0;
	1273: instructionOdd = 32'h0;
	1274: instructionOdd = 32'h0;
	1275: instructionOdd = 32'h0;
	1276: instructionOdd = 32'h0;
	1277: instructionOdd = 32'h0;
	1278: instructionOdd = 32'h0;
	1279: instructionOdd = 32'h0;
	1280: instructionOdd = 32'h0;
	1281: instructionOdd = 32'h0;
	1282: instructionOdd = 32'h0;
	1283: instructionOdd = 32'h0;
	1284: instructionOdd = 32'h0;
	1285: instructionOdd = 32'h0;
	1286: instructionOdd = 32'h0;
	1287: instructionOdd = 32'h0;
	1288: instructionOdd = 32'h0;
	1289: instructionOdd = 32'h0;
	1290: instructionOdd = 32'h0;
	1291: instructionOdd = 32'h0;
	1292: instructionOdd = 32'h0;
	1293: instructionOdd = 32'h0;
	1294: instructionOdd = 32'h0;
	1295: instructionOdd = 32'h0;
	1296: instructionOdd = 32'h0;
	1297: instructionOdd = 32'h0;
	1298: instructionOdd = 32'h0;
	1299: instructionOdd = 32'h0;
	1300: instructionOdd = 32'h0;
	1301: instructionOdd = 32'h0;
	1302: instructionOdd = 32'h0;
	1303: instructionOdd = 32'h0;
	1304: instructionOdd = 32'h0;
	1305: instructionOdd = 32'h0;
	1306: instructionOdd = 32'h0;
	1307: instructionOdd = 32'h0;
	1308: instructionOdd = 32'h0;
	1309: instructionOdd = 32'h0;
	1310: instructionOdd = 32'h0;
	1311: instructionOdd = 32'h0;
	1312: instructionOdd = 32'h0;
	1313: instructionOdd = 32'h0;
	1314: instructionOdd = 32'h0;
	1315: instructionOdd = 32'h0;
	1316: instructionOdd = 32'h0;
	1317: instructionOdd = 32'h0;
	1318: instructionOdd = 32'h0;
	1319: instructionOdd = 32'h0;
	1320: instructionOdd = 32'h0;
	1321: instructionOdd = 32'h0;
	1322: instructionOdd = 32'h0;
	1323: instructionOdd = 32'h0;
	1324: instructionOdd = 32'h0;
	1325: instructionOdd = 32'h0;
	1326: instructionOdd = 32'h0;
	1327: instructionOdd = 32'h0;
	1328: instructionOdd = 32'h0;
	1329: instructionOdd = 32'h0;
	1330: instructionOdd = 32'h0;
	1331: instructionOdd = 32'h0;
	1332: instructionOdd = 32'h0;
	1333: instructionOdd = 32'h0;
	1334: instructionOdd = 32'h0;
	1335: instructionOdd = 32'h0;
	1336: instructionOdd = 32'h0;
	1337: instructionOdd = 32'h0;
	1338: instructionOdd = 32'h0;
	1339: instructionOdd = 32'h0;
	1340: instructionOdd = 32'h0;
	1341: instructionOdd = 32'h0;
	1342: instructionOdd = 32'h0;
	1343: instructionOdd = 32'h0;
	1344: instructionOdd = 32'h0;
	1345: instructionOdd = 32'h0;
	1346: instructionOdd = 32'h0;
	1347: instructionOdd = 32'h0;
	1348: instructionOdd = 32'h0;
	1349: instructionOdd = 32'h0;
	1350: instructionOdd = 32'h0;
	1351: instructionOdd = 32'h0;
	1352: instructionOdd = 32'h0;
	1353: instructionOdd = 32'h0;
	1354: instructionOdd = 32'h0;
	1355: instructionOdd = 32'h0;
	1356: instructionOdd = 32'h0;
	1357: instructionOdd = 32'h0;
	1358: instructionOdd = 32'h0;
	1359: instructionOdd = 32'h0;
	1360: instructionOdd = 32'h0;
	1361: instructionOdd = 32'h0;
	1362: instructionOdd = 32'h0;
	1363: instructionOdd = 32'h0;
	1364: instructionOdd = 32'h0;
	1365: instructionOdd = 32'h0;
	1366: instructionOdd = 32'h0;
	1367: instructionOdd = 32'h0;
	1368: instructionOdd = 32'h0;
	1369: instructionOdd = 32'h0;
	1370: instructionOdd = 32'h0;
	1371: instructionOdd = 32'h0;
	1372: instructionOdd = 32'h0;
	1373: instructionOdd = 32'h0;
	1374: instructionOdd = 32'h0;
	1375: instructionOdd = 32'h0;
	1376: instructionOdd = 32'h0;
	1377: instructionOdd = 32'h0;
	1378: instructionOdd = 32'h0;
	1379: instructionOdd = 32'h0;
	1380: instructionOdd = 32'h0;
	1381: instructionOdd = 32'h0;
	1382: instructionOdd = 32'h0;
	1383: instructionOdd = 32'h0;
	1384: instructionOdd = 32'h0;
	1385: instructionOdd = 32'h0;
	1386: instructionOdd = 32'h0;
	1387: instructionOdd = 32'h0;
	1388: instructionOdd = 32'h0;
	1389: instructionOdd = 32'h0;
	1390: instructionOdd = 32'h0;
	1391: instructionOdd = 32'h0;
	1392: instructionOdd = 32'h0;
	1393: instructionOdd = 32'h0;
	1394: instructionOdd = 32'h0;
	1395: instructionOdd = 32'h0;
	1396: instructionOdd = 32'h0;
	1397: instructionOdd = 32'h0;
	1398: instructionOdd = 32'h0;
	1399: instructionOdd = 32'h0;
	1400: instructionOdd = 32'h0;
	1401: instructionOdd = 32'h0;
	1402: instructionOdd = 32'h0;
	1403: instructionOdd = 32'h0;
	1404: instructionOdd = 32'h0;
	1405: instructionOdd = 32'h0;
	1406: instructionOdd = 32'h0;
	1407: instructionOdd = 32'h0;
	1408: instructionOdd = 32'h0;
	1409: instructionOdd = 32'h0;
	1410: instructionOdd = 32'h0;
	1411: instructionOdd = 32'h0;
	1412: instructionOdd = 32'h0;
	1413: instructionOdd = 32'h0;
	1414: instructionOdd = 32'h0;
	1415: instructionOdd = 32'h0;
	1416: instructionOdd = 32'h0;
	1417: instructionOdd = 32'h0;
	1418: instructionOdd = 32'h0;
	1419: instructionOdd = 32'h0;
	1420: instructionOdd = 32'h0;
	1421: instructionOdd = 32'h0;
	1422: instructionOdd = 32'h0;
	1423: instructionOdd = 32'h0;
	1424: instructionOdd = 32'h0;
	1425: instructionOdd = 32'h0;
	1426: instructionOdd = 32'h0;
	1427: instructionOdd = 32'h0;
	1428: instructionOdd = 32'h0;
	1429: instructionOdd = 32'h0;
	1430: instructionOdd = 32'h0;
	1431: instructionOdd = 32'h0;
	1432: instructionOdd = 32'h0;
	1433: instructionOdd = 32'h0;
	1434: instructionOdd = 32'h0;
	1435: instructionOdd = 32'h0;
	1436: instructionOdd = 32'h0;
	1437: instructionOdd = 32'h0;
	1438: instructionOdd = 32'h0;
	1439: instructionOdd = 32'h0;
	1440: instructionOdd = 32'h0;
	1441: instructionOdd = 32'h0;
	1442: instructionOdd = 32'h0;
	1443: instructionOdd = 32'h0;
	1444: instructionOdd = 32'h0;
	1445: instructionOdd = 32'h0;
	1446: instructionOdd = 32'h0;
	1447: instructionOdd = 32'h0;
	1448: instructionOdd = 32'h0;
	1449: instructionOdd = 32'h0;
	1450: instructionOdd = 32'h0;
	1451: instructionOdd = 32'h0;
	1452: instructionOdd = 32'h0;
	1453: instructionOdd = 32'h0;
	1454: instructionOdd = 32'h0;
	1455: instructionOdd = 32'h0;
	1456: instructionOdd = 32'h0;
	1457: instructionOdd = 32'h0;
	1458: instructionOdd = 32'h0;
	1459: instructionOdd = 32'h0;
	1460: instructionOdd = 32'h0;
	1461: instructionOdd = 32'h0;
	1462: instructionOdd = 32'h0;
	1463: instructionOdd = 32'h0;
	1464: instructionOdd = 32'h0;
	1465: instructionOdd = 32'h0;
	1466: instructionOdd = 32'h0;
	1467: instructionOdd = 32'h0;
	1468: instructionOdd = 32'h0;
	1469: instructionOdd = 32'h0;
	1470: instructionOdd = 32'h0;
	1471: instructionOdd = 32'h0;
	1472: instructionOdd = 32'h0;
	1473: instructionOdd = 32'h0;
	1474: instructionOdd = 32'h0;
	1475: instructionOdd = 32'h0;
	1476: instructionOdd = 32'h0;
	1477: instructionOdd = 32'h0;
	1478: instructionOdd = 32'h0;
	1479: instructionOdd = 32'h0;
	1480: instructionOdd = 32'h0;
	1481: instructionOdd = 32'h0;
	1482: instructionOdd = 32'h0;
	1483: instructionOdd = 32'h0;
	1484: instructionOdd = 32'h0;
	1485: instructionOdd = 32'h0;
	1486: instructionOdd = 32'h0;
	1487: instructionOdd = 32'h0;
	1488: instructionOdd = 32'h0;
	1489: instructionOdd = 32'h0;
	1490: instructionOdd = 32'h0;
	1491: instructionOdd = 32'h0;
	1492: instructionOdd = 32'h0;
	1493: instructionOdd = 32'h0;
	1494: instructionOdd = 32'h0;
	1495: instructionOdd = 32'h0;
	1496: instructionOdd = 32'h0;
	1497: instructionOdd = 32'h0;
	1498: instructionOdd = 32'h0;
	1499: instructionOdd = 32'h0;
	1500: instructionOdd = 32'h0;
	1501: instructionOdd = 32'h0;
	1502: instructionOdd = 32'h0;
	1503: instructionOdd = 32'h0;
	1504: instructionOdd = 32'h0;
	1505: instructionOdd = 32'h0;
	1506: instructionOdd = 32'h0;
	1507: instructionOdd = 32'h0;
	1508: instructionOdd = 32'h0;
	1509: instructionOdd = 32'h0;
	1510: instructionOdd = 32'h0;
	1511: instructionOdd = 32'h0;
	1512: instructionOdd = 32'h0;
	1513: instructionOdd = 32'h0;
	1514: instructionOdd = 32'h0;
	1515: instructionOdd = 32'h0;
	1516: instructionOdd = 32'h0;
	1517: instructionOdd = 32'h0;
	1518: instructionOdd = 32'h0;
	1519: instructionOdd = 32'h0;
	1520: instructionOdd = 32'h0;
	1521: instructionOdd = 32'h0;
	1522: instructionOdd = 32'h0;
	1523: instructionOdd = 32'h0;
	1524: instructionOdd = 32'h0;
	1525: instructionOdd = 32'h0;
	1526: instructionOdd = 32'h0;
	1527: instructionOdd = 32'h0;
	1528: instructionOdd = 32'h0;
	1529: instructionOdd = 32'h0;
	1530: instructionOdd = 32'h0;
	1531: instructionOdd = 32'h0;
	1532: instructionOdd = 32'h0;
	1533: instructionOdd = 32'h0;
	1534: instructionOdd = 32'h0;
	1535: instructionOdd = 32'h0;
	1536: instructionOdd = 32'h0;
	1537: instructionOdd = 32'h0;
	1538: instructionOdd = 32'h0;
	1539: instructionOdd = 32'h0;
	1540: instructionOdd = 32'h0;
	1541: instructionOdd = 32'h0;
	1542: instructionOdd = 32'h0;
	1543: instructionOdd = 32'h0;
	1544: instructionOdd = 32'h0;
	1545: instructionOdd = 32'h0;
	1546: instructionOdd = 32'h0;
	1547: instructionOdd = 32'h0;
	1548: instructionOdd = 32'h0;
	1549: instructionOdd = 32'h0;
	1550: instructionOdd = 32'h0;
	1551: instructionOdd = 32'h0;
	1552: instructionOdd = 32'h0;
	1553: instructionOdd = 32'h0;
	1554: instructionOdd = 32'h0;
	1555: instructionOdd = 32'h0;
	1556: instructionOdd = 32'h0;
	1557: instructionOdd = 32'h0;
	1558: instructionOdd = 32'h0;
	1559: instructionOdd = 32'h0;
	1560: instructionOdd = 32'h0;
	1561: instructionOdd = 32'h0;
	1562: instructionOdd = 32'h0;
	1563: instructionOdd = 32'h0;
	1564: instructionOdd = 32'h0;
	1565: instructionOdd = 32'h0;
	1566: instructionOdd = 32'h0;
	1567: instructionOdd = 32'h0;
	1568: instructionOdd = 32'h0;
	1569: instructionOdd = 32'h0;
	1570: instructionOdd = 32'h0;
	1571: instructionOdd = 32'h0;
	1572: instructionOdd = 32'h0;
	1573: instructionOdd = 32'h0;
	1574: instructionOdd = 32'h0;
	1575: instructionOdd = 32'h0;
	1576: instructionOdd = 32'h0;
	1577: instructionOdd = 32'h0;
	1578: instructionOdd = 32'h0;
	1579: instructionOdd = 32'h0;
	1580: instructionOdd = 32'h0;
	1581: instructionOdd = 32'h0;
	1582: instructionOdd = 32'h0;
	1583: instructionOdd = 32'h0;
	1584: instructionOdd = 32'h0;
	1585: instructionOdd = 32'h0;
	1586: instructionOdd = 32'h0;
	1587: instructionOdd = 32'h0;
	1588: instructionOdd = 32'h0;
	1589: instructionOdd = 32'h0;
	1590: instructionOdd = 32'h0;
	1591: instructionOdd = 32'h0;
	1592: instructionOdd = 32'h0;
	1593: instructionOdd = 32'h0;
	1594: instructionOdd = 32'h0;
	1595: instructionOdd = 32'h0;
	1596: instructionOdd = 32'h0;
	1597: instructionOdd = 32'h0;
	1598: instructionOdd = 32'h0;
	1599: instructionOdd = 32'h0;
	1600: instructionOdd = 32'h0;
	1601: instructionOdd = 32'h0;
	1602: instructionOdd = 32'h0;
	1603: instructionOdd = 32'h0;
	1604: instructionOdd = 32'h0;
	1605: instructionOdd = 32'h0;
	1606: instructionOdd = 32'h0;
	1607: instructionOdd = 32'h0;
	1608: instructionOdd = 32'h0;
	1609: instructionOdd = 32'h0;
	1610: instructionOdd = 32'h0;
	1611: instructionOdd = 32'h0;
	1612: instructionOdd = 32'h0;
	1613: instructionOdd = 32'h0;
	1614: instructionOdd = 32'h0;
	1615: instructionOdd = 32'h0;
	1616: instructionOdd = 32'h0;
	1617: instructionOdd = 32'h0;
	1618: instructionOdd = 32'h0;
	1619: instructionOdd = 32'h0;
	1620: instructionOdd = 32'h0;
	1621: instructionOdd = 32'h0;
	1622: instructionOdd = 32'h0;
	1623: instructionOdd = 32'h0;
	1624: instructionOdd = 32'h0;
	1625: instructionOdd = 32'h0;
	1626: instructionOdd = 32'h0;
	1627: instructionOdd = 32'h0;
	1628: instructionOdd = 32'h0;
	1629: instructionOdd = 32'h0;
	1630: instructionOdd = 32'h0;
	1631: instructionOdd = 32'h0;
	1632: instructionOdd = 32'h0;
	1633: instructionOdd = 32'h0;
	1634: instructionOdd = 32'h0;
	1635: instructionOdd = 32'h0;
	1636: instructionOdd = 32'h0;
	1637: instructionOdd = 32'h0;
	1638: instructionOdd = 32'h0;
	1639: instructionOdd = 32'h0;
	1640: instructionOdd = 32'h0;
	1641: instructionOdd = 32'h0;
	1642: instructionOdd = 32'h0;
	1643: instructionOdd = 32'h0;
	1644: instructionOdd = 32'h0;
	1645: instructionOdd = 32'h0;
	1646: instructionOdd = 32'h0;
	1647: instructionOdd = 32'h0;
	1648: instructionOdd = 32'h0;
	1649: instructionOdd = 32'h0;
	1650: instructionOdd = 32'h0;
	1651: instructionOdd = 32'h0;
	1652: instructionOdd = 32'h0;
	1653: instructionOdd = 32'h0;
	1654: instructionOdd = 32'h0;
	1655: instructionOdd = 32'h0;
	1656: instructionOdd = 32'h0;
	1657: instructionOdd = 32'h0;
	1658: instructionOdd = 32'h0;
	1659: instructionOdd = 32'h0;
	1660: instructionOdd = 32'h0;
	1661: instructionOdd = 32'h0;
	1662: instructionOdd = 32'h0;
	1663: instructionOdd = 32'h0;
	1664: instructionOdd = 32'h0;
	1665: instructionOdd = 32'h0;
	1666: instructionOdd = 32'h0;
	1667: instructionOdd = 32'h0;
	1668: instructionOdd = 32'h0;
	1669: instructionOdd = 32'h0;
	1670: instructionOdd = 32'h0;
	1671: instructionOdd = 32'h0;
	1672: instructionOdd = 32'h0;
	1673: instructionOdd = 32'h0;
	1674: instructionOdd = 32'h0;
	1675: instructionOdd = 32'h0;
	1676: instructionOdd = 32'h0;
	1677: instructionOdd = 32'h0;
	1678: instructionOdd = 32'h0;
	1679: instructionOdd = 32'h0;
	1680: instructionOdd = 32'h0;
	1681: instructionOdd = 32'h0;
	1682: instructionOdd = 32'h0;
	1683: instructionOdd = 32'h0;
	1684: instructionOdd = 32'h0;
	1685: instructionOdd = 32'h0;
	1686: instructionOdd = 32'h0;
	1687: instructionOdd = 32'h0;
	1688: instructionOdd = 32'h0;
	1689: instructionOdd = 32'h0;
	1690: instructionOdd = 32'h0;
	1691: instructionOdd = 32'h0;
	1692: instructionOdd = 32'h0;
	1693: instructionOdd = 32'h0;
	1694: instructionOdd = 32'h0;
	1695: instructionOdd = 32'h0;
	1696: instructionOdd = 32'h0;
	1697: instructionOdd = 32'h0;
	1698: instructionOdd = 32'h0;
	1699: instructionOdd = 32'h0;
	1700: instructionOdd = 32'h0;
	1701: instructionOdd = 32'h0;
	1702: instructionOdd = 32'h0;
	1703: instructionOdd = 32'h0;
	1704: instructionOdd = 32'h0;
	1705: instructionOdd = 32'h0;
	1706: instructionOdd = 32'h0;
	1707: instructionOdd = 32'h0;
	1708: instructionOdd = 32'h0;
	1709: instructionOdd = 32'h0;
	1710: instructionOdd = 32'h0;
	1711: instructionOdd = 32'h0;
	1712: instructionOdd = 32'h0;
	1713: instructionOdd = 32'h0;
	1714: instructionOdd = 32'h0;
	1715: instructionOdd = 32'h0;
	1716: instructionOdd = 32'h0;
	1717: instructionOdd = 32'h0;
	1718: instructionOdd = 32'h0;
	1719: instructionOdd = 32'h0;
	1720: instructionOdd = 32'h0;
	1721: instructionOdd = 32'h0;
	1722: instructionOdd = 32'h0;
	1723: instructionOdd = 32'h0;
	1724: instructionOdd = 32'h0;
	1725: instructionOdd = 32'h0;
	1726: instructionOdd = 32'h0;
	1727: instructionOdd = 32'h0;
	1728: instructionOdd = 32'h0;
	1729: instructionOdd = 32'h0;
	1730: instructionOdd = 32'h0;
	1731: instructionOdd = 32'h0;
	1732: instructionOdd = 32'h0;
	1733: instructionOdd = 32'h0;
	1734: instructionOdd = 32'h0;
	1735: instructionOdd = 32'h0;
	1736: instructionOdd = 32'h0;
	1737: instructionOdd = 32'h0;
	1738: instructionOdd = 32'h0;
	1739: instructionOdd = 32'h0;
	1740: instructionOdd = 32'h0;
	1741: instructionOdd = 32'h0;
	1742: instructionOdd = 32'h0;
	1743: instructionOdd = 32'h0;
	1744: instructionOdd = 32'h0;
	1745: instructionOdd = 32'h0;
	1746: instructionOdd = 32'h0;
	1747: instructionOdd = 32'h0;
	1748: instructionOdd = 32'h0;
	1749: instructionOdd = 32'h0;
	1750: instructionOdd = 32'h0;
	1751: instructionOdd = 32'h0;
	1752: instructionOdd = 32'h0;
	1753: instructionOdd = 32'h0;
	1754: instructionOdd = 32'h0;
	1755: instructionOdd = 32'h0;
	1756: instructionOdd = 32'h0;
	1757: instructionOdd = 32'h0;
	1758: instructionOdd = 32'h0;
	1759: instructionOdd = 32'h0;
	1760: instructionOdd = 32'h0;
	1761: instructionOdd = 32'h0;
	1762: instructionOdd = 32'h0;
	1763: instructionOdd = 32'h0;
	1764: instructionOdd = 32'h0;
	1765: instructionOdd = 32'h0;
	1766: instructionOdd = 32'h0;
	1767: instructionOdd = 32'h0;
	1768: instructionOdd = 32'h0;
	1769: instructionOdd = 32'h0;
	1770: instructionOdd = 32'h0;
	1771: instructionOdd = 32'h0;
	1772: instructionOdd = 32'h0;
	1773: instructionOdd = 32'h0;
	1774: instructionOdd = 32'h0;
	1775: instructionOdd = 32'h0;
	1776: instructionOdd = 32'h0;
	1777: instructionOdd = 32'h0;
	1778: instructionOdd = 32'h0;
	1779: instructionOdd = 32'h0;
	1780: instructionOdd = 32'h0;
	1781: instructionOdd = 32'h0;
	1782: instructionOdd = 32'h0;
	1783: instructionOdd = 32'h0;
	1784: instructionOdd = 32'h0;
	1785: instructionOdd = 32'h0;
	1786: instructionOdd = 32'h0;
	1787: instructionOdd = 32'h0;
	1788: instructionOdd = 32'h0;
	1789: instructionOdd = 32'h0;
	1790: instructionOdd = 32'h0;
	1791: instructionOdd = 32'h0;
	1792: instructionOdd = 32'h0;
	1793: instructionOdd = 32'h0;
	1794: instructionOdd = 32'h0;
	1795: instructionOdd = 32'h0;
	1796: instructionOdd = 32'h0;
	1797: instructionOdd = 32'h0;
	1798: instructionOdd = 32'h0;
	1799: instructionOdd = 32'h0;
	1800: instructionOdd = 32'h0;
	1801: instructionOdd = 32'h0;
	1802: instructionOdd = 32'h0;
	1803: instructionOdd = 32'h0;
	1804: instructionOdd = 32'h0;
	1805: instructionOdd = 32'h0;
	1806: instructionOdd = 32'h0;
	1807: instructionOdd = 32'h0;
	1808: instructionOdd = 32'h0;
	1809: instructionOdd = 32'h0;
	1810: instructionOdd = 32'h0;
	1811: instructionOdd = 32'h0;
	1812: instructionOdd = 32'h0;
	1813: instructionOdd = 32'h0;
	1814: instructionOdd = 32'h0;
	1815: instructionOdd = 32'h0;
	1816: instructionOdd = 32'h0;
	1817: instructionOdd = 32'h0;
	1818: instructionOdd = 32'h0;
	1819: instructionOdd = 32'h0;
	1820: instructionOdd = 32'h0;
	1821: instructionOdd = 32'h0;
	1822: instructionOdd = 32'h0;
	1823: instructionOdd = 32'h0;
	1824: instructionOdd = 32'h0;
	1825: instructionOdd = 32'h0;
	1826: instructionOdd = 32'h0;
	1827: instructionOdd = 32'h0;
	1828: instructionOdd = 32'h0;
	1829: instructionOdd = 32'h0;
	1830: instructionOdd = 32'h0;
	1831: instructionOdd = 32'h0;
	1832: instructionOdd = 32'h0;
	1833: instructionOdd = 32'h0;
	1834: instructionOdd = 32'h0;
	1835: instructionOdd = 32'h0;
	1836: instructionOdd = 32'h0;
	1837: instructionOdd = 32'h0;
	1838: instructionOdd = 32'h0;
	1839: instructionOdd = 32'h0;
	1840: instructionOdd = 32'h0;
	1841: instructionOdd = 32'h0;
	1842: instructionOdd = 32'h0;
	1843: instructionOdd = 32'h0;
	1844: instructionOdd = 32'h0;
	1845: instructionOdd = 32'h0;
	1846: instructionOdd = 32'h0;
	1847: instructionOdd = 32'h0;
	1848: instructionOdd = 32'h0;
	1849: instructionOdd = 32'h0;
	1850: instructionOdd = 32'h0;
	1851: instructionOdd = 32'h0;
	1852: instructionOdd = 32'h0;
	1853: instructionOdd = 32'h0;
	1854: instructionOdd = 32'h0;
	1855: instructionOdd = 32'h0;
	1856: instructionOdd = 32'h0;
	1857: instructionOdd = 32'h0;
	1858: instructionOdd = 32'h0;
	1859: instructionOdd = 32'h0;
	1860: instructionOdd = 32'h0;
	1861: instructionOdd = 32'h0;
	1862: instructionOdd = 32'h0;
	1863: instructionOdd = 32'h0;
	1864: instructionOdd = 32'h0;
	1865: instructionOdd = 32'h0;
	1866: instructionOdd = 32'h0;
	1867: instructionOdd = 32'h0;
	1868: instructionOdd = 32'h0;
	1869: instructionOdd = 32'h0;
	1870: instructionOdd = 32'h0;
	1871: instructionOdd = 32'h0;
	1872: instructionOdd = 32'h0;
	1873: instructionOdd = 32'h0;
	1874: instructionOdd = 32'h0;
	1875: instructionOdd = 32'h0;
	1876: instructionOdd = 32'h0;
	1877: instructionOdd = 32'h0;
	1878: instructionOdd = 32'h0;
	1879: instructionOdd = 32'h0;
	1880: instructionOdd = 32'h0;
	1881: instructionOdd = 32'h0;
	1882: instructionOdd = 32'h0;
	1883: instructionOdd = 32'h0;
	1884: instructionOdd = 32'h0;
	1885: instructionOdd = 32'h0;
	1886: instructionOdd = 32'h0;
	1887: instructionOdd = 32'h0;
	1888: instructionOdd = 32'h0;
	1889: instructionOdd = 32'h0;
	1890: instructionOdd = 32'h0;
	1891: instructionOdd = 32'h0;
	1892: instructionOdd = 32'h0;
	1893: instructionOdd = 32'h0;
	1894: instructionOdd = 32'h0;
	1895: instructionOdd = 32'h0;
	1896: instructionOdd = 32'h0;
	1897: instructionOdd = 32'h0;
	1898: instructionOdd = 32'h0;
	1899: instructionOdd = 32'h0;
	1900: instructionOdd = 32'h0;
	1901: instructionOdd = 32'h0;
	1902: instructionOdd = 32'h0;
	1903: instructionOdd = 32'h0;
	1904: instructionOdd = 32'h0;
	1905: instructionOdd = 32'h0;
	1906: instructionOdd = 32'h0;
	1907: instructionOdd = 32'h0;
	1908: instructionOdd = 32'h0;
	1909: instructionOdd = 32'h0;
	1910: instructionOdd = 32'h0;
	1911: instructionOdd = 32'h0;
	1912: instructionOdd = 32'h0;
	1913: instructionOdd = 32'h0;
	1914: instructionOdd = 32'h0;
	1915: instructionOdd = 32'h0;
	1916: instructionOdd = 32'h0;
	1917: instructionOdd = 32'h0;
	1918: instructionOdd = 32'h0;
	1919: instructionOdd = 32'h0;
	1920: instructionOdd = 32'h0;
	1921: instructionOdd = 32'h0;
	1922: instructionOdd = 32'h0;
	1923: instructionOdd = 32'h0;
	1924: instructionOdd = 32'h0;
	1925: instructionOdd = 32'h0;
	1926: instructionOdd = 32'h0;
	1927: instructionOdd = 32'h0;
	1928: instructionOdd = 32'h0;
	1929: instructionOdd = 32'h0;
	1930: instructionOdd = 32'h0;
	1931: instructionOdd = 32'h0;
	1932: instructionOdd = 32'h0;
	1933: instructionOdd = 32'h0;
	1934: instructionOdd = 32'h0;
	1935: instructionOdd = 32'h0;
	1936: instructionOdd = 32'h0;
	1937: instructionOdd = 32'h0;
	1938: instructionOdd = 32'h0;
	1939: instructionOdd = 32'h0;
	1940: instructionOdd = 32'h0;
	1941: instructionOdd = 32'h0;
	1942: instructionOdd = 32'h0;
	1943: instructionOdd = 32'h0;
	1944: instructionOdd = 32'h0;
	1945: instructionOdd = 32'h0;
	1946: instructionOdd = 32'h0;
	1947: instructionOdd = 32'h0;
	1948: instructionOdd = 32'h0;
	1949: instructionOdd = 32'h0;
	1950: instructionOdd = 32'h0;
	1951: instructionOdd = 32'h0;
	1952: instructionOdd = 32'h0;
	1953: instructionOdd = 32'h0;
	1954: instructionOdd = 32'h0;
	1955: instructionOdd = 32'h0;
	1956: instructionOdd = 32'h0;
	1957: instructionOdd = 32'h0;
	1958: instructionOdd = 32'h0;
	1959: instructionOdd = 32'h0;
	1960: instructionOdd = 32'h0;
	1961: instructionOdd = 32'h0;
	1962: instructionOdd = 32'h0;
	1963: instructionOdd = 32'h0;
	1964: instructionOdd = 32'h0;
	1965: instructionOdd = 32'h0;
	1966: instructionOdd = 32'h0;
	1967: instructionOdd = 32'h0;
	1968: instructionOdd = 32'h0;
	1969: instructionOdd = 32'h0;
	1970: instructionOdd = 32'h0;
	1971: instructionOdd = 32'h0;
	1972: instructionOdd = 32'h0;
	1973: instructionOdd = 32'h0;
	1974: instructionOdd = 32'h0;
	1975: instructionOdd = 32'h0;
	1976: instructionOdd = 32'h0;
	1977: instructionOdd = 32'h0;
	1978: instructionOdd = 32'h0;
	1979: instructionOdd = 32'h0;
	1980: instructionOdd = 32'h0;
	1981: instructionOdd = 32'h0;
	1982: instructionOdd = 32'h0;
	1983: instructionOdd = 32'h0;
	1984: instructionOdd = 32'h0;
	1985: instructionOdd = 32'h0;
	1986: instructionOdd = 32'h0;
	1987: instructionOdd = 32'h0;
	1988: instructionOdd = 32'h0;
	1989: instructionOdd = 32'h0;
	1990: instructionOdd = 32'h0;
	1991: instructionOdd = 32'h0;
	1992: instructionOdd = 32'h0;
	1993: instructionOdd = 32'h0;
	1994: instructionOdd = 32'h0;
	1995: instructionOdd = 32'h0;
	1996: instructionOdd = 32'h0;
	1997: instructionOdd = 32'h0;
	1998: instructionOdd = 32'h0;
	1999: instructionOdd = 32'h0;
	2000: instructionOdd = 32'h0;
	2001: instructionOdd = 32'h0;
	2002: instructionOdd = 32'h0;
	2003: instructionOdd = 32'h0;
	2004: instructionOdd = 32'h0;
	2005: instructionOdd = 32'h0;
	2006: instructionOdd = 32'h0;
	2007: instructionOdd = 32'h0;
	2008: instructionOdd = 32'h0;
	2009: instructionOdd = 32'h0;
	2010: instructionOdd = 32'h0;
	2011: instructionOdd = 32'h0;
	2012: instructionOdd = 32'h0;
	2013: instructionOdd = 32'h0;
	2014: instructionOdd = 32'h0;
	2015: instructionOdd = 32'h0;
	2016: instructionOdd = 32'h0;
	2017: instructionOdd = 32'h0;
	2018: instructionOdd = 32'h0;
	2019: instructionOdd = 32'h0;
	2020: instructionOdd = 32'h0;
	2021: instructionOdd = 32'h0;
	2022: instructionOdd = 32'h0;
	2023: instructionOdd = 32'h0;
	2024: instructionOdd = 32'h0;
	2025: instructionOdd = 32'h0;
	2026: instructionOdd = 32'h0;
	2027: instructionOdd = 32'h0;
	2028: instructionOdd = 32'h0;
	2029: instructionOdd = 32'h0;
	2030: instructionOdd = 32'h0;
	2031: instructionOdd = 32'h0;
	2032: instructionOdd = 32'h0;
	2033: instructionOdd = 32'h0;
	2034: instructionOdd = 32'h0;
	2035: instructionOdd = 32'h0;
	2036: instructionOdd = 32'h0;
	2037: instructionOdd = 32'h0;
	2038: instructionOdd = 32'h0;
	2039: instructionOdd = 32'h0;
	2040: instructionOdd = 32'h0;
	2041: instructionOdd = 32'h0;
	2042: instructionOdd = 32'h0;
	2043: instructionOdd = 32'h0;
	2044: instructionOdd = 32'h0;
	2045: instructionOdd = 32'h0;
	2046: instructionOdd = 32'h0;
	2047: instructionOdd = 32'h0;

    default: begin
        instructionOdd = 32'bx;
        `ifndef SYNTHESIS
            // synthesis translate_off
            instructionOdd = {1{$random}};
            // synthesis translate_on
        `endif
    end
endcase
        
endmodule
